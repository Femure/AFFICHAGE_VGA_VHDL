LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY memory_rom IS
	PORT (
		RST : IN STD_LOGIC;
		HCOUNT, VCOUNT : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		RED, GREEN, BLUE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END memory_rom;

ARCHITECTURE rtl OF memory_rom IS

	TYPE data_Array IS ARRAY (0 TO 60160) OF STD_LOGIC_VECTOR(11 DOWNTO 0);

	-- Initialisation des données
	CONSTANT XMAX : INTEGER := 600;
	CONSTANT YMAX : INTEGER := 315;

	CONSTANT data_vector : data_Array := (
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"101010000111",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"101010000111",
		"011101000011",
		"011101000011",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111011101111",
		"111011101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111011101111",
		"110111101111",
		"110111101111",
		"110111101111",
		"111011101111",
		"110111101111",
		"110111101111",
		"111011101111",
		"111011101111",
		"111111101110",
		"111111101110",
		"111111101101",
		"111111011101",
		"111111011101",
		"111111101101",
		"111111101101",
		"111111101101",
		"111111011101",
		"111111011101",
		"111111011101",
		"111111011101",
		"111111101101",
		"111111101101",
		"111111101101",
		"111111011100",
		"101010000111",
		"100001000011",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101000011",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011101111010",
		"010001001001",
		"010001001010",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001001011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001001011",
		"010001001011",
		"010001001011",
		"010101001010",
		"011001000111",
		"011001000101",
		"011001000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000010",
		"100001000011",
		"100001000011",
		"100001000011",
		"011101000011",
		"011101000010",
		"011101000010",
		"100001000011",
		"011100110010",
		"100000110010",
		"100101000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001011",
		"011001000111",
		"011101000100",
		"011101000010",
		"011101000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100100110001",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011100",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001011",
		"011101000111",
		"011100110100",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001011",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"001101011100",
		"001101011100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010101001011",
		"011101000111",
		"011100110100",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011101",
		"001101001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101001100",
		"010001011101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010101001011",
		"011101000111",
		"011101000100",
		"100001000011",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010101001011",
		"011001000111",
		"011101000100",
		"011101000011",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001011",
		"011001010111",
		"011101000100",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001011",
		"011001010111",
		"011101000100",
		"011101000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001100",
		"001101011101",
		"001101001101",
		"010001001011",
		"011001000111",
		"011101000011",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001011",
		"011001000111",
		"011101000011",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001011",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100001000001",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001111100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010101011100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110010",
		"100001000011",
		"100001000011",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011001101011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001010011",
		"011000110010",
		"011101000011",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001011",
		"111011001100",
		"110111001101",
		"110111001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"110011001111",
		"101111001111",
		"010101101100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011100110010",
		"100101100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"100001100101",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000011",
		"011001000100",
		"011001000110",
		"010101001000",
		"010001011010",
		"010101011010",
		"010101011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001001010",
		"010001001010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001001010",
		"010001001010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001001010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001011010",
		"010001001010",
		"010001001010",
		"010101011010",
		"010001011011",
		"010001011010",
		"010001001010",
		"010001011011",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"011101000010",
		"110110111010",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111110",
		"111111111111",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"011101000011",
		"011101000100",
		"011001000110",
		"010101001010",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001011100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001011100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001011100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001011",
		"010001011100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110110111010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000010",
		"110110111010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000101",
		"010101001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001110",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000011",
		"110110111010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000101",
		"010101001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"011101000011",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000101",
		"010101001010",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"011101000011",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100101000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000101",
		"010101001010",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001011101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"011101000011",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110011",
		"011101000110",
		"010001001011",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001010",
		"011001000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110001",
		"011101000010",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110011",
		"011101000110",
		"010001001011",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"011101000111",
		"011101000100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110010",
		"011101000011",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010101001011",
		"011101000111",
		"011101000100",
		"011100110010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"011101000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100000110010",
		"011101000011",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"001101001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001010",
		"011101000111",
		"011101000100",
		"100001000011",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110001",
		"100000110001",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"100001000001",
		"100000110001",
		"100001000010",
		"011101000011",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011100110011",
		"011001000101",
		"010001001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001011101",
		"001101001101",
		"001101001100",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"001101011100",
		"001101011100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"001101001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001011",
		"011101000111",
		"011100110011",
		"011100110010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000001",
		"011101000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"011100110010",
		"110010111010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101001100",
		"001101001100",
		"001101011101",
		"001101001101",
		"010001011101",
		"010001011100",
		"010001011100",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011100",
		"010001011100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011100",
		"010001011100",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001011",
		"011101000111",
		"011100110100",
		"100001000011",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100000110010",
		"100001000010",
		"011101000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000101",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101001100",
		"001101001100",
		"010001011101",
		"001101001101",
		"001101001100",
		"010001011100",
		"010001011101",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011101",
		"010001001101",
		"001101001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001010",
		"011001000111",
		"011101000100",
		"011101000011",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110110111010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000101",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011100",
		"010001011011",
		"010001011010",
		"010001011001",
		"010001011010",
		"010001011011",
		"010001001011",
		"010001001011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010101011010",
		"010101011010",
		"010101011010",
		"010001011011",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010101001011",
		"011001011000",
		"011001000100",
		"011101000011",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000011",
		"011101000011",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000011",
		"110010111010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000011",
		"011101000110",
		"010101011010",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010101011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010101011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001011100",
		"010001001010",
		"011001101010",
		"011001100111",
		"011001100110",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001100111",
		"011001101001",
		"010101011011",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010101011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010101011101",
		"010001001101",
		"010001011101",
		"010101001011",
		"011101011000",
		"100001100110",
		"011101010101",
		"100001100100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010101",
		"100001010101",
		"011101010100",
		"011101010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001100101",
		"011101010100",
		"100001010100",
		"100001010100",
		"100001010100",
		"100001100101",
		"110010111011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001011",
		"010101011010",
		"101110111101",
		"110111011011",
		"111011101010",
		"111011101010",
		"111011011010",
		"111011011010",
		"111011101010",
		"111011101010",
		"111011101010",
		"111011101010",
		"111011101010",
		"111011101010",
		"111011101010",
		"110111101001",
		"111011101001",
		"111011101010",
		"110111011101",
		"010001011010",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011011",
		"101010011100",
		"111111101111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001011",
		"111011101000",
		"111011100110",
		"111011100110",
		"111111100101",
		"111111100101",
		"111111100101",
		"111011100101",
		"111011100101",
		"111011100101",
		"111011100101",
		"111011100110",
		"111011100110",
		"111011100101",
		"111011100101",
		"111011100110",
		"111011101010",
		"010101011001",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011011",
		"101010011100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111011100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111011101000",
		"010101011001",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011011",
		"100110011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111011101000",
		"010101011001",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011011",
		"100110011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111110011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111011101000",
		"010101011001",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011100",
		"100110011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111011101000",
		"010101011001",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011011",
		"100110011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001011011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111011101000",
		"010101011001",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011011",
		"100110011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011011",
		"010101010111",
		"110011001010",
		"111011100110",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111011101000",
		"010001011000",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011011",
		"100110011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011011",
		"010101010111",
		"110011001010",
		"111011100110",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111011101000",
		"010001011000",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"101010011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101011100",
		"001101001100",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001011100",
		"010001011100",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111101000",
		"010101011001",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011100",
		"001101011100",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"101010011100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011101",
		"001101011100",
		"001101001100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011100",
		"010001011100",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101001100",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111011101000",
		"010101011001",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"001101011100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"100110011100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001010",
		"111011100110",
		"111111110100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111110011",
		"111111110011",
		"111111110100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111101000",
		"010101011001",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011100",
		"001101001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"001101011100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"100110011100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101011101",
		"001101011101",
		"001101011101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101010111",
		"110011001010",
		"111011100110",
		"111011100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111011100100",
		"111011100100",
		"111011100100",
		"111011100100",
		"111011100100",
		"111011100100",
		"111011100100",
		"111111100100",
		"111111100100",
		"111011101000",
		"010101011001",
		"001101011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101011100",
		"001101001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011100",
		"010001011100",
		"001101011100",
		"001101011101",
		"001101001100",
		"010001001101",
		"010001001101",
		"010001011011",
		"100110101100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001110",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001010",
		"010101010111",
		"110011001010",
		"111011100110",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111011101000",
		"010101011001",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"100110101100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001011101",
		"001101001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001010",
		"010101010111",
		"110011001010",
		"111011100111",
		"111011100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100101",
		"111111100101",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111011100100",
		"111111100100",
		"111111100100",
		"111011101000",
		"010101011001",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001011",
		"100110101100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"001101011100",
		"001101001100",
		"001101001100",
		"010001011100",
		"010001011011",
		"010001001011",
		"010001011011",
		"010001001011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001011100",
		"010001001100",
		"010001011101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001011",
		"010101011000",
		"110011001011",
		"111011101000",
		"111011100101",
		"111111100101",
		"111111100101",
		"111111100100",
		"111111100101",
		"111111100101",
		"111111100101",
		"111111100101",
		"111111100101",
		"111111100101",
		"111111100101",
		"111011100101",
		"111111100101",
		"111111100101",
		"111011101001",
		"010101011001",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001100",
		"010101001101",
		"010101001101",
		"010001001100",
		"010101001100",
		"010101001100",
		"010101001010",
		"101010011100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011100",
		"010001011100",
		"010001001100",
		"010001011100",
		"010101101010",
		"011001101001",
		"011001101001",
		"011001111001",
		"011001111001",
		"011001111001",
		"011001101001",
		"011001101001",
		"011001111001",
		"011001111001",
		"011001111001",
		"011001101001",
		"011001101001",
		"011001101010",
		"011001101001",
		"011001101001",
		"011001101010",
		"010101101011",
		"010001011100",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001001",
		"101110111100",
		"110011001001",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011001000",
		"110011001000",
		"110011001000",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011000111",
		"110011001010",
		"010101011010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"011100111001",
		"011100111000",
		"011100111001",
		"011100111001",
		"011100111001",
		"011100111010",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111000",
		"100001001001",
		"100000111000",
		"100000111001",
		"100000111000",
		"100000111000",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111000",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111000",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111001",
		"100000111000",
		"101101111001",
		"111111001100",
		"111110111100",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111110111011",
		"111111001100",
		"111111011110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010101001010",
		"101010101010",
		"111011101010",
		"111011101001",
		"111011101000",
		"111011101000",
		"111011100111",
		"111011100111",
		"111011100111",
		"111011100111",
		"111011101000",
		"111011101000",
		"111011101000",
		"111011101000",
		"111011101000",
		"111011101000",
		"111011101001",
		"110111011011",
		"100010001001",
		"010001001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001011011",
		"010001011010",
		"010001011000",
		"010001011000",
		"010001011001",
		"010001011001",
		"010001011001",
		"010001011000",
		"010001011000",
		"010001011000",
		"010001011001",
		"010001011001",
		"010001011000",
		"010001011000",
		"010001011001",
		"010001011000",
		"010001011000",
		"010001011001",
		"010001011100",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"011100111010",
		"101000010101",
		"110000000011",
		"110000010010",
		"110000010010",
		"110000000010",
		"110000000011",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110100010011",
		"110000000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110000000010",
		"110000010010",
		"110100010011",
		"110000010010",
		"110000000010",
		"110000010010",
		"110100000010",
		"110000010010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110000010011",
		"110000000011",
		"110000000011",
		"110100000011",
		"110100010010",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110000010001",
		"101000100010",
		"111010011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"010101001001",
		"101010101000",
		"111011100111",
		"111011100101",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111011100101",
		"111011101000",
		"100010000111",
		"010001001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101011101",
		"001101001101",
		"001101011100",
		"010001011100",
		"010001011100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"001101011100",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001011101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000011",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111110001000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001001",
		"101010100111",
		"111011100110",
		"111011100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100101",
		"111011101000",
		"100010000111",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001011",
		"100000111001",
		"110000000011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"111110001000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010101001010",
		"101010100111",
		"111011100110",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111011101000",
		"100010000111",
		"010001001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"001101011100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110001000",
		"111111101111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001110",
		"010101001010",
		"101010100111",
		"111011100110",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111011101000",
		"100010000111",
		"010001001010",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"100000111001",
		"110000000011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010101001010",
		"101010101000",
		"111011100110",
		"111111100101",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001011010",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"100000111001",
		"110000000011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010101001001",
		"101010101000",
		"111011100111",
		"111111100101",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001011010",
		"001101001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000011",
		"011101000110",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"010001001100",
		"010001001100",
		"010101001001",
		"101010101000",
		"111011100111",
		"111111100101",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100110",
		"111011101000",
		"100010000111",
		"010001011010",
		"001101011101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000101",
		"010101001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011001",
		"101010101000",
		"111011100111",
		"111111100101",
		"111111100011",
		"111111110011",
		"111111110011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001011010",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010000",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000101",
		"010101001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011001",
		"101010101000",
		"111111100111",
		"111111100101",
		"111111100011",
		"111011110011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001011010",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010000",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000101",
		"010101001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011010",
		"101010101000",
		"111111100111",
		"111111100101",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001001010",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000101",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001011010",
		"101010101000",
		"111111100110",
		"111111100101",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100101",
		"111111011000",
		"100010000111",
		"010101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011001000101",
		"010101001010",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"001101001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001011001",
		"101010100111",
		"111111100110",
		"111111100101",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000101",
		"010101001010",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011001",
		"101010101000",
		"111011100111",
		"111111100101",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100100",
		"111111100100",
		"111111100011",
		"111111100101",
		"111011101000",
		"100010000111",
		"010001001010",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"011001000110",
		"010101001010",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011001",
		"101010101000",
		"111011100111",
		"111011100101",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111111100011",
		"111011100011",
		"111011100100",
		"111111100100",
		"111111100011",
		"111111100011",
		"111111110011",
		"111011100101",
		"110111101000",
		"100010000111",
		"010001001010",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111110001000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011100110011",
		"011101000110",
		"010101001001",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001001100",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001011",
		"010001001011",
		"010001001011",
		"010001001100",
		"010001001100",
		"010101011100",
		"010001001011",
		"010001001100",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001011",
		"010001011011",
		"010101011000",
		"101010101001",
		"111011101001",
		"111011101000",
		"111011100111",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100110",
		"111011100111",
		"111011101010",
		"100010001000",
		"011001001000",
		"011001001010",
		"011001001011",
		"010101001011",
		"010101001010",
		"010101001010",
		"010101001010",
		"010101001010",
		"011001001010",
		"011001001011",
		"011001001011",
		"011001001010",
		"011001001011",
		"011001001011",
		"011001001010",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001010",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"010101001011",
		"010101001011",
		"011001001011",
		"011001001011",
		"011001001010",
		"010101001011",
		"010001001101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111110000111",
		"111111101110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101010011",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000011",
		"011101010101",
		"100010001011",
		"011110001100",
		"011101111100",
		"100010001100",
		"011101111100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011110001100",
		"011101111011",
		"100010001011",
		"100110011010",
		"101010101010",
		"101110111011",
		"101010111001",
		"101110111001",
		"101110111001",
		"101110111010",
		"101110111010",
		"101110111010",
		"101110111010",
		"101110111010",
		"101110111010",
		"101110111010",
		"101110101001",
		"101110111010",
		"101110111010",
		"101110101010",
		"101001111000",
		"101000110110",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000111000",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"101000110111",
		"100100111000",
		"011001011100",
		"010001011110",
		"010001011101",
		"010101011101",
		"010101011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010001011101",
		"010101011101",
		"010101001100",
		"100001001001",
		"110100010011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111000010001",
		"111101100101",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011010",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011010",
		"111110011001",
		"111110011001",
		"111110011001",
		"111110011001",
		"111111101110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101100101",
		"111111101111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111011101111",
		"100010001011",
		"010101011000",
		"010001011000",
		"010101011000",
		"010101011000",
		"010101011000",
		"010101011001",
		"010101011001",
		"010101001001",
		"010101001001",
		"010101001000",
		"010101001000",
		"010101011001",
		"010001011000",
		"010001011000",
		"010101011000",
		"011101001000",
		"100000110110",
		"101000010011",
		"110000000011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"101100010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010100",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000000011",
		"110000000011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"110000010011",
		"101000010101",
		"011001001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001011101",
		"010001001101",
		"010001001101",
		"010101001100",
		"100000111001",
		"110100010010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"110100000000",
		"110100010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"101100100010",
		"111010101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001011011",
		"010001001011",
		"010001011011",
		"010001011011",
		"010001011011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010101001100",
		"010101001100",
		"010001001100",
		"010001001100",
		"010001001011",
		"010001001010",
		"011100111001",
		"101000100111",
		"110100010011",
		"111100000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111100000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"101100010011",
		"011101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110100000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011110001101",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001110",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001100",
		"011100111010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011101001010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001011",
		"011100111010",
		"101000100110",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010010",
		"011101001010",
		"001101001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100101100101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010011101",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011101",
		"010001001101",
		"001101011101",
		"010001001011",
		"011101001010",
		"101000100111",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011101001010",
		"010001001101",
		"001101001100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001100100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001100",
		"001101001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001011100",
		"010001001100",
		"010001001100",
		"001101001100",
		"001101011100",
		"010001001011",
		"011100111010",
		"101000100111",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011100111010",
		"010001001100",
		"010001001100",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001100",
		"010001011011",
		"010001011100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001011100",
		"010001001011",
		"011100111010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011100111010",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001011",
		"011100111010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011101001010",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001011",
		"011101001010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011101001010",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001001011",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001011101",
		"010001001011",
		"011001001010",
		"100100100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011101001010",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101011101",
		"001101011100",
		"010001011100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010101001100",
		"100000111001",
		"110000000011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001001011",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"010001011101",
		"010001001011",
		"011001001010",
		"100100100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011100111010",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"001101011100",
		"001101011100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"100000111001",
		"110100000011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001011011",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010101001100",
		"011100111010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011100111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001011",
		"100000111000",
		"110100000011",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"100001100100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001101",
		"010001011011",
		"010001001100",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010101001100",
		"011100111010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011100111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001011",
		"100000111000",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001100101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001100",
		"010001011011",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"011100111010",
		"101000100111",
		"110100000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010011",
		"011101001010",
		"001101011101",
		"001101001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010101001100",
		"100000111000",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000011",
		"100001100101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100010001100",
		"010101001010",
		"010001001011",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010101001100",
		"010101001100",
		"010001001101",
		"010101001011",
		"011100111001",
		"101000100110",
		"110100000010",
		"111100000000",
		"111000000000",
		"111000000000",
		"111100000001",
		"111100000001",
		"111100000001",
		"111100000001",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111000000001",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010010",
		"011101001001",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010101001011",
		"100000111000",
		"110000010010",
		"111100000000",
		"111000000000",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000011",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011001000011",
		"011101100101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100110001100",
		"011001001010",
		"011001001011",
		"011001001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001010",
		"100000111000",
		"101000100110",
		"110000010011",
		"110100000010",
		"110100010001",
		"110100000001",
		"110100000001",
		"111000000010",
		"111000000010",
		"111000000010",
		"110100000010",
		"110100000010",
		"110100000001",
		"110100010001",
		"110100000001",
		"110100000001",
		"110100000010",
		"111000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000010",
		"100000111000",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"011001001011",
		"011001001011",
		"011001001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"011001001011",
		"100000111000",
		"101100010011",
		"110100000001",
		"110100000010",
		"111000000010",
		"111000000001",
		"110100000001",
		"110100000001",
		"110100000001",
		"110100000001",
		"110100000001",
		"110100000010",
		"110100000010",
		"111000000001",
		"111000000010",
		"110100000010",
		"111000000010",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"101110000110",
		"101110000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111011001100",
		"110110011001",
		"111010011001",
		"111010011001",
		"111010011001",
		"111010011001",
		"111010011001",
		"111010011001",
		"111110011001",
		"111110011001",
		"111110011001",
		"111010011001",
		"111010011001",
		"111110011001",
		"111010011001",
		"111010011001",
		"111010001010",
		"101001011000",
		"100000100111",
		"100000101000",
		"100000101000",
		"100000101000",
		"100000101000",
		"100000101000",
		"100000101000",
		"100000100111",
		"100000100111",
		"100000101000",
		"100000101000",
		"100000101000",
		"100000100111",
		"100000101000",
		"100000100111",
		"100100100110",
		"101000100110",
		"101000100101",
		"101000100101",
		"101000100101",
		"101000100101",
		"101100010101",
		"101100010101",
		"101100010101",
		"101100010101",
		"101100010101",
		"101100010101",
		"101000100101",
		"101000100101",
		"101000100101",
		"101000100101",
		"101100100101",
		"110000010100",
		"111000000010",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"101000100110",
		"100000100111",
		"100100100111",
		"100100100111",
		"100100100111",
		"100000100111",
		"100000101000",
		"100000101000",
		"100000100111",
		"100000100111",
		"100000100111",
		"100100101000",
		"100000100111",
		"100000100111",
		"100000110111",
		"100000110111",
		"100000100111",
		"100100100111",
		"101000100101",
		"101000100101",
		"101100010110",
		"101100010110",
		"101100010101",
		"101100100100",
		"101100100101",
		"101000100101",
		"101100100101",
		"101100100101",
		"101000100101",
		"101100100101",
		"101100010101",
		"101100010101",
		"101100010101",
		"110000010101",
		"111000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100101100101",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"110110001000",
		"101100100010",
		"110000010001",
		"110100000001",
		"110100000001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100000000",
		"110100010001",
		"110100000000",
		"110100010001",
		"110100010010",
		"110100000010",
		"110100010011",
		"110100000011",
		"110100000011",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110000010010",
		"110000010010",
		"110000000010",
		"110000010011",
		"101100010100",
		"100100110111",
		"011100111001",
		"011001001010",
		"010101001010",
		"010101001011",
		"011000111010",
		"011100111010",
		"011100111010",
		"011000111010",
		"011000111010",
		"011000111010",
		"011000111011",
		"011000111011",
		"011000111010",
		"011000111010",
		"011100111001",
		"100100101000",
		"110000010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000010",
		"110100000011",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000010",
		"110100000011",
		"110100000011",
		"110100000010",
		"110100010010",
		"110100000010",
		"110100000010",
		"110100010010",
		"110100010010",
		"110100010001",
		"110100010010",
		"110000010011",
		"101100010101",
		"100000111000",
		"011001001010",
		"011000111011",
		"011000111011",
		"011001001010",
		"011001001010",
		"011000111010",
		"011000111010",
		"011000111010",
		"011000111010",
		"011001001011",
		"011001001011",
		"011001001010",
		"011001001010",
		"011000111010",
		"100000111000",
		"101100100101",
		"110000010010",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111010000111",
		"110000010001",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000110111",
		"011001001010",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010101001100",
		"011100111001",
		"110000010101",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"101100010100",
		"011001001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101011101",
		"010001001100",
		"010001001100",
		"011001001010",
		"101000110111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111010001000",
		"110100000001",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000110111",
		"011001001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"001101011100",
		"001101011100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001100",
		"010001001100",
		"011100111001",
		"110000010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"101100010101",
		"011001001010",
		"001101011101",
		"010001001101",
		"010001001101",
		"001101011100",
		"001101011100",
		"001101011100",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"011001001011",
		"101000110111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010100",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111001111000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000100111",
		"011001001011",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001011100",
		"001101011101",
		"001101011101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101001101",
		"010001001100",
		"011100111010",
		"110000010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000001",
		"111000000001",
		"101100010101",
		"011000111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101001100",
		"001101011101",
		"010001001100",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011000111011",
		"101000100111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001100101",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111010000111",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000100111",
		"010101001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001110",
		"001101001110",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"011001001010",
		"101100100100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010100",
		"011100111001",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"001101011100",
		"010001001101",
		"011001001011",
		"101000100111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111010000111",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000000011",
		"101000100111",
		"010101001011",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001110",
		"010001001110",
		"010001001110",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"011000111010",
		"101100010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010100",
		"011100111001",
		"010001001100",
		"010001001100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011100",
		"001101011100",
		"001101011101",
		"011001001011",
		"101000110111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111010000111",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000100111",
		"011001001011",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001110",
		"010001001110",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"010001001100",
		"011100111010",
		"101100010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010100",
		"011100111001",
		"010001001100",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011100",
		"010001011100",
		"010001001101",
		"011001001011",
		"101000110111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111010101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111010000111",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000100111",
		"011001001011",
		"010001001101",
		"010001011100",
		"010001011100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011100",
		"010001001100",
		"011100111010",
		"101100010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"101100010100",
		"011100111010",
		"010001001101",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001011100",
		"010001001100",
		"010001001101",
		"011001001011",
		"101000110111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111010101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111010001000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000000011",
		"101000100111",
		"011001001011",
		"010001001101",
		"010001001100",
		"010001001100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"011100111010",
		"101100010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"101100010100",
		"011100111010",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"010001001100",
		"010001001100",
		"010001001101",
		"011001001011",
		"101000100111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111010001000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000000011",
		"101000100111",
		"011001001011",
		"010001001101",
		"010001001100",
		"010001001100",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011100111010",
		"101100010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"101100010101",
		"011100111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"011001001011",
		"101000100111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111010001000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000110111",
		"010101001011",
		"010001011101",
		"010001001100",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011000111010",
		"101100010100",
		"111000000001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000001",
		"101100010101",
		"011000111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001100",
		"010001001100",
		"011001001011",
		"101000110111",
		"110000010011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111010001000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010011",
		"101000110111",
		"011001001011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011000111010",
		"101100010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"101100010100",
		"011000111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"010001001101",
		"011001001011",
		"101000110111",
		"110000010011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111001111000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000100111",
		"011000111011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101011101",
		"001101011101",
		"001101001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011000111010",
		"110000010100",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010100",
		"011000111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101001101",
		"001101011101",
		"001101011101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011000111011",
		"101000100111",
		"110000010011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"011101000010",
		"100001010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111010001000",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"101000100111",
		"011000111011",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011100",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011100111010",
		"110000010100",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010100",
		"011100111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"001101011101",
		"001101011100",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011000111011",
		"101000100111",
		"110000010011",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111110101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101010100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111001110111",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010011",
		"100100100111",
		"011001001010",
		"010001001100",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"001101011101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"011100111010",
		"110000010100",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000001",
		"110000010100",
		"011100111010",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001101",
		"010001001100",
		"011001001010",
		"100100100111",
		"110000010011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111110101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000011",
		"011101010101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111101111",
		"111111111111",
		"111111111111",
		"111111101111",
		"111111101111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111101101",
		"111101110111",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000010000",
		"110100000000",
		"110100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000010000",
		"111000000000",
		"110100010001",
		"101100100011",
		"100100110110",
		"011001001001",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010101001010",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"011100111001",
		"101100100100",
		"110100010001",
		"110100000001",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000010000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110100000001",
		"110100010001",
		"101100100100",
		"011100111000",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001011",
		"010101001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"010001001010",
		"011001001001",
		"100100110110",
		"101100100011",
		"110100010000",
		"111000000000",
		"111000010000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110100000000",
		"111000000000",
		"111000010000",
		"111000010001",
		"110100000001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010001",
		"110100010000",
		"110100010000",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100000000",
		"110100000001",
		"110100000000",
		"101100010001",
		"111110101010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110011000",
		"101110101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111011101",
		"111010000111",
		"111101110111",
		"111101110110",
		"111101110111",
		"111101110111",
		"111101100111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101110111",
		"111101000100",
		"111100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111100000000",
		"111000010000",
		"111101010011",
		"111101110101",
		"111101100101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110100",
		"111101110101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"110101110110",
		"110010001000",
		"101010001010",
		"100110001010",
		"100110001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"100110001011",
		"101010001001",
		"110101110110",
		"111101110101",
		"111101100101",
		"111101100101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111001110101",
		"111101110101",
		"111101110101",
		"111101100101",
		"111101110101",
		"111101110101",
		"111101100101",
		"111101100101",
		"111101110101",
		"111101110101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101100101",
		"111101110101",
		"111001110101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111001110101",
		"110101110110",
		"101010001001",
		"100110001011",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"101010001010",
		"100110001010",
		"101010001010",
		"110010001000",
		"111001110110",
		"111101100101",
		"111101100100",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101100101",
		"111101110101",
		"111101110101",
		"111101110101",
		"111001110110",
		"111110000111",
		"111001110111",
		"111001110111",
		"111001110111",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111010001000",
		"111001111000",
		"111001111000",
		"111010001000",
		"111010001000",
		"111010001000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111001111000",
		"111010001000",
		"111010001000",
		"111010001000",
		"111001111000",
		"111010001000",
		"111001111000",
		"111001110111",
		"111001110111",
		"111001111000",
		"111001111000",
		"111001110111",
		"111001110111",
		"111010000111",
		"111010001000",
		"111010001000",
		"111010001000",
		"111001111000",
		"110110001001",
		"111011011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"101100100010",
		"110100000000",
		"110100010000",
		"110100010001",
		"110100010001",
		"110100000001",
		"110100010001",
		"110100010001",
		"110100010000",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100000001",
		"110100010001",
		"110100010001",
		"111000010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010000",
		"111101110101",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111010",
		"111010111011",
		"110110111011",
		"111010111011",
		"111010111011",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"110110111010",
		"111010111010",
		"110110111011",
		"110110111011",
		"111010111010",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111010111010",
		"110110111011",
		"110110111011",
		"111010111010",
		"110110111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111011",
		"111010111011",
		"110110111011",
		"111010111011",
		"111110111010",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111010",
		"111111101101",
		"111111101110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000001",
		"111000000000",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111010",
		"111010111010",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111010",
		"111010111010",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111011001001",
		"110111001010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111011001000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001001",
		"111011001001",
		"110111001010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111001110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111011001000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"110111001010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111011001001",
		"110111001010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111011001001",
		"110111001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111101110101",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111011001001",
		"110111001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111101110101",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111011001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111011001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"110111001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111011001001",
		"110111001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111001",
		"111010111000",
		"111011001001",
		"111011001001",
		"110111001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111011001001",
		"111011001001",
		"111011001001",
		"111010111000",
		"111010111000",
		"111111001001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111011001001",
		"111010111000",
		"110111001001",
		"110111001010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"110100000000",
		"111101110101",
		"111110111001",
		"111110111001",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111111001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111011001001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111011001001",
		"111011001000",
		"111011001001",
		"110111001010",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000010000",
		"110100000000",
		"110100010001",
		"110100000001",
		"111000000001",
		"111000000001",
		"111000000001",
		"110100000001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110100010001",
		"110000010001",
		"110101110110",
		"111110111001",
		"111010111001",
		"111011001001",
		"111011001001",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111011001001",
		"111011001001",
		"111011001001",
		"111011001001",
		"110110111001",
		"111111001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111011001000",
		"111011001001",
		"110111001001",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000000000",
		"100000000000",
		"011100000000",
		"100000000000",
		"100000000000",
		"100000000000",
		"100000000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011100000000",
		"011000000000",
		"011100110010",
		"011101000011",
		"011001000011",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011101010011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001010011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001010011",
		"011001000010",
		"011001010011",
		"011001000011",
		"011001000011",
		"011001000010",
		"011101010011",
		"110110111000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111011001001",
		"111010111000",
		"110010100111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"101010000111",
		"100110001000",
		"110111001100",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"101000000000",
		"010000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"000100000000",
		"000100000000",
		"000100000000",
		"000100000000",
		"000100000000",
		"001000000000",
		"001000000000",
		"000100000000",
		"000100000000",
		"001000000000",
		"000100000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"101110010110",
		"011101000010",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100000001",
		"100100000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010111001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"110010010110",
		"011100110010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100001000001",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100100000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"110010010110",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100000110010",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101001",
		"111011001001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"110010000101",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010000",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111000",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111000",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111011001001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"110010000110",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100000000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111011001001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"110010000110",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010000",
		"100100000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111011001001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"110010000110",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010000",
		"100000000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111110111001",
		"110010000110",
		"100001000001",
		"100001000010",
		"100000110001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010001",
		"100100000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"000000000000",
		"110010101001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111011111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111110111011",
		"110000010001",
		"111100000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"100100000000",
		"001000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111111001001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"110010000110",
		"011101000001",
		"011100110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111111110",
		"111111111110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101111",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111111111110",
		"111110101001",
		"110000100010",
		"110100000000",
		"110100000000",
		"110100010000",
		"110100010000",
		"110100000000",
		"110100000000",
		"111000000000",
		"110100000000",
		"110100000000",
		"110100000000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"101100010000",
		"100000000000",
		"001100000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"000100000000",
		"001000000000",
		"110010101000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111111001001",
		"111111001001",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"110010000110",
		"100001000010",
		"011101000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"011100110001",
		"011101000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000001",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111011100",
		"101101010101",
		"111001010101",
		"111101010101",
		"111101000100",
		"111101000100",
		"111001010100",
		"111001010100",
		"111001010100",
		"111001010100",
		"111001010100",
		"111001010101",
		"111001010100",
		"111001010100",
		"111001010100",
		"111001010100",
		"111001000100",
		"111101010101",
		"111110000111",
		"111110000111",
		"111110000110",
		"111010000110",
		"111110010110",
		"111110010110",
		"111110000110",
		"111110000110",
		"111110000111",
		"111110000111",
		"111110000110",
		"111110010110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110010110",
		"110110010110",
		"101110000110",
		"101110010111",
		"101010010111",
		"101110010111",
		"101110000111",
		"101110000111",
		"101110000111",
		"101110000111",
		"101110010111",
		"101110010111",
		"101010010111",
		"101010010111",
		"101110010111",
		"101110010111",
		"101110010110",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110010110",
		"101110010111",
		"101110010110",
		"101110010111",
		"101110010110",
		"101110010111",
		"101110010110",
		"101110010111",
		"101110010110",
		"101110010111",
		"101010000110",
		"101010000111",
		"101010000111",
		"101010011000",
		"101010011000",
		"010101000011",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000010000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"000100000000",
		"100001110110",
		"101010010111",
		"101010010111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101010000111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110010111",
		"101110000111",
		"101110000110",
		"111010111001",
		"111011001001",
		"111011001001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111111001000",
		"111111001000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010101000",
		"101001110100",
		"101001110100",
		"101001110100",
		"101101110100",
		"101101110100",
		"101101110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001100100",
		"101001110100",
		"101001110100",
		"110010000110",
		"110110010111",
		"110110100111",
		"110110010111",
		"110110100111",
		"110110010111",
		"110110010111",
		"110110010111",
		"110110010111",
		"110110010111",
		"110110010111",
		"110110010111",
		"110110010111",
		"110110100111",
		"110110010111",
		"110110010111",
		"110110010111",
		"101101110101",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101000010",
		"100101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101000010",
		"100101000010",
		"100101000010",
		"100101000010",
		"100001000011",
		"100001000011",
		"110110101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"101000100001",
		"110100010001",
		"111000000001",
		"111000000000",
		"111000000000",
		"110100000000",
		"110100010000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110100000000",
		"110100000000",
		"111000000000",
		"111000000000",
		"111000000001",
		"111000100010",
		"111110101000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110110111",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"110110111010",
		"110111001010",
		"010101000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"000100000000",
		"101110010111",
		"111011001010",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001010",
		"111010111001",
		"111011001001",
		"111111001001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"110110100111",
		"100001000010",
		"100001000010",
		"011101000001",
		"100001000001",
		"100001000001",
		"011100110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"101101110101",
		"111110111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001011",
		"101100010001",
		"111000000001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000110010",
		"111110101000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111111001000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111011001001",
		"111011001001",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111001",
		"111011001001",
		"111011001010",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"101110010111",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001000",
		"111010111000",
		"111010111001",
		"111111001001",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110100111",
		"011101000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"011101000001",
		"101101110101",
		"111010111000",
		"111110111001",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111001",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000001",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"101100010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000110010",
		"111110101000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111111001001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001001",
		"110110111001",
		"011001000010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"101110010111",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111111001000",
		"111111001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"110110100111",
		"011101000001",
		"100001000010",
		"011100110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"101101110101",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"110010000110",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000100010",
		"111110101000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111110111001",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110011000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111001",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000110",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000100010",
		"111110101000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110011000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000100010",
		"111110101000",
		"111110111000",
		"111010111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000110010",
		"111110101000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000110010",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111010111000",
		"111010111001",
		"111010111010",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000110010",
		"111110111000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111010111000",
		"111010111001",
		"111010111010",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000110010",
		"111110111000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000100010",
		"111110101000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111011001001",
		"111011001001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000100010",
		"111110111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111011001001",
		"111010111000",
		"111010111000",
		"111111001001",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111111001000",
		"111010111000",
		"111011001001",
		"010101000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111111001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"011100110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000110010",
		"111110101000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111011001001",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110010111",
		"111010111001",
		"111010111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000110010",
		"111110101000",
		"111010111000",
		"111111001000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111111001000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111010111001",
		"111011001010",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"101110011000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111011001001",
		"111011001001",
		"111011001001",
		"111011001001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000001",
		"011101000001",
		"011100110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111100110010",
		"111110010111",
		"111110111000",
		"111110111000",
		"111110101000",
		"111110101000",
		"111110111000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110111000",
		"111110101000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"110110111000",
		"011001000010",
		"000100000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"101010010111",
		"111011001010",
		"111011001010",
		"111011001010",
		"111011001010",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"110110111001",
		"110110111001",
		"110110111001",
		"111011001001",
		"110110111001",
		"111111001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"110110010111",
		"100001000010",
		"100001000001",
		"011101000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100000110001",
		"100000110001",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111101000011",
		"111101010011",
		"111101010011",
		"111101010011",
		"111101010100",
		"111101010100",
		"111101010011",
		"111101010011",
		"111101010011",
		"111101010011",
		"111101010011",
		"111101010100",
		"111101010100",
		"111101010100",
		"111101010100",
		"111101010100",
		"111001010100",
		"111110000110",
		"111110111000",
		"111110111000",
		"111110111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111111001000",
		"111010111001",
		"101110010110",
		"100101110101",
		"100001110101",
		"100001110101",
		"100001110101",
		"100101110101",
		"100101110101",
		"100101110101",
		"100101110101",
		"100101110101",
		"100101110101",
		"100001110101",
		"100101110101",
		"100101110101",
		"100101110101",
		"100101110101",
		"100001100101",
		"011101100100",
		"011001010011",
		"011001010011",
		"011001010100",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001010011",
		"011001010100",
		"011001010011",
		"011001000011",
		"011001010011",
		"011101010011",
		"110110111000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"110010000110",
		"101101110101",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110100000000",
		"110000010000",
		"111101100100",
		"111110101000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"110110111001",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001010",
		"111010111001",
		"111010111000",
		"111010111001",
		"111011001001",
		"110110111001",
		"010000110001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111111001001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100000110001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110100010000",
		"111101100100",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111001",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111111001001",
		"111010111001",
		"111010111001",
		"111011001010",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111111001001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111101100100",
		"111110101000",
		"111110111000",
		"111010111000",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111111001001",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111011001001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"110110010111",
		"011101000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100101",
		"111110101000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"011101000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111010111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100001000001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100101",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111001",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100100",
		"111110111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111011001000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"110010000110",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000001",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100100",
		"111110101000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"101101110101",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110010000110",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100100",
		"111110101000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000001",
		"101101110101",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110010000110",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000001",
		"100000110001",
		"100000110001",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100100",
		"111110101000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000001",
		"101101110101",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100000110010",
		"100001000010",
		"011101000011",
		"110010101010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101100100",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000001",
		"101101110101",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000011",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101100101",
		"111110111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111011001001",
		"111010111000",
		"111011001001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000110001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000001",
		"011101000001",
		"101101110101",
		"111110111001",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000001",
		"100000110001",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100000110001",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101100101",
		"111110101000",
		"111010111000",
		"111010111000",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111011001001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"010000110001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"101101110101",
		"111110111001",
		"111010111000",
		"111111001001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110010000101",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110001",
		"100000110001",
		"100000110001",
		"100000110001",
		"100000110001",
		"100000110001",
		"100001000010",
		"100000110001",
		"100001000001",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111101100100",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111111001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111001",
		"111010111001",
		"010000110010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"101101110101",
		"111110111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"110010000101",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011100110001",
		"100001000010",
		"100001000010",
		"011101000010",
		"110010101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010010",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111101010100",
		"111110101000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111011001001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"111011001010",
		"111011001001",
		"111010111001",
		"111010111001",
		"111111001001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111110111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111001",
		"110110010111",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000001",
		"101101110101",
		"111110111001",
		"111110111001",
		"111110111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"101110000110",
		"011101000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"110010101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"101100010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000010000",
		"111101010100",
		"111110100111",
		"111110111000",
		"111110101000",
		"111110111000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110100111",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110111001",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"111010111010",
		"110110111010",
		"110110111010",
		"110110111010",
		"110110111010",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000110010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"110110010111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"101101110101",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010111001",
		"101110000110",
		"011101000011",
		"011001000010",
		"011101000011",
		"011101000011",
		"011101000011",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000010",
		"011101000011",
		"011101000011",
		"011001000011",
		"011001000011",
		"011101000011",
		"011101000010",
		"011101010011",
		"110010101001",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000100010",
		"111100010001",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111000000000",
		"111100110010",
		"111101010011",
		"111001010011",
		"111001000011",
		"111001000011",
		"111001000011",
		"111001010011",
		"110101010011",
		"110101010011",
		"111001010011",
		"111001000011",
		"111001000011",
		"111001000011",
		"111001010011",
		"111101010011",
		"111001000011",
		"110101010100",
		"110110011000",
		"111011011011",
		"111011011011",
		"111011011011",
		"111111001011",
		"111111001100",
		"111011011100",
		"111011011100",
		"111011011011",
		"111011001011",
		"111011011011",
		"111011011011",
		"111011011100",
		"111011011100",
		"111011011100",
		"111011011011",
		"111111011011",
		"111010111001",
		"111011001001",
		"111011001001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111111001001",
		"111010111001",
		"111011001001",
		"111111001001",
		"111011001001",
		"010000110010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110110111001",
		"111011001001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010101000",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001110100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001110100",
		"101101110100",
		"101001100100",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100101010011",
		"101101110100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001110100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001100100",
		"101001110101",
		"101110010111",
		"110110111010",
		"110110111010",
		"110110111011",
		"110110111011",
		"110110111011",
		"110110111010",
		"110110111010",
		"110110111010",
		"110110111010",
		"110110111011",
		"110110111011",
		"110111001011",
		"110110111010",
		"110110111010",
		"110110111010",
		"110110111010",
		"111011011101",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111000010000",
		"110100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000010000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110100000000",
		"110000010001",
		"111010011000",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"111111111101",
		"110110111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000110010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"110110100111",
		"100001000010",
		"011101000001",
		"011101000001",
		"011101000001",
		"011101000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011100110001",
		"011100110001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"101110011000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"110110111001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"010000110010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110101000",
		"011101000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110001",
		"100001000010",
		"100001000010",
		"100000110001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100000110001",
		"100000110001",
		"100000110001",
		"100001000010",
		"100001000010",
		"011101000010",
		"101110011000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"110110111010",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"001100100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"011101000010",
		"101110011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"001100100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"011101000010",
		"101110011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"001100100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"110110100111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"011101000010",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"110110100111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"011101000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"011101000011",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010000",
		"111010001000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"110110100111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"011101000010",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010011000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"110110111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"011101000010",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111010111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"010000100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"011101000010",
		"101110011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111010001001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111010111001",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111011001001",
		"001100100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"110110100111",
		"100001000001",
		"100001000001",
		"100001000010",
		"100000110001",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"011101000010",
		"101110011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111110",
		"110110111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111011001010",
		"010000100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111001",
		"110110100111",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"011101000001",
		"011101000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100000110001",
		"100001000001",
		"100001000001",
		"100001000010",
		"011101000010",
		"101110101000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111011",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111001",
		"010000100010",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000100000000",
		"110010101001",
		"111010111001",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"110110100111",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"011101000001",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100000110001",
		"100000110001",
		"100000110010",
		"100001000001",
		"100001000001",
		"100001000010",
		"011101000010",
		"101110101000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010000",
		"111010011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111011001001",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111001",
		"010000110001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010101000",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"110110101000",
		"011100110001",
		"011101000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111110111100",
		"101100010001",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010000",
		"111010011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110010111010",
		"111010111001",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111111001001",
		"111111001001",
		"111110111000",
		"111010111001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111010101000",
		"011101000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100000110010",
		"100000110010",
		"100001000010",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"011101000010",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"110000010010",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000010001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"110110111010",
		"111011001001",
		"111011001001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111010111001",
		"111010111000",
		"111010111000",
		"111011001001",
		"010000100001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010111001",
		"111010111001",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010100111",
		"011100110001",
		"100001000001",
		"100001000001",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100000110010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000010",
		"100001000001",
		"100000110001",
		"100001000010",
		"100001000010",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100001000001",
		"100000110001",
		"100000110010",
		"011101000010",
		"101110011001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111001100",
		"101100100010",
		"110100010000",
		"110100000000",
		"110100000000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100000000",
		"110100000000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100000000",
		"111000010000",
		"111100000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000010001",
		"111110001000",
		"111111011110",
		"111111101110",
		"111111101110",
		"111111111110",
		"111111111110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111111101110",
		"111110101001",
		"111110101000",
		"111110101000",
		"111110101001",
		"111110101001",
		"111110111000",
		"111110111000",
		"111110101000",
		"111110101000",
		"111110111000",
		"111110101000",
		"111110111000",
		"111110101000",
		"111110111000",
		"111110101000",
		"111110101000",
		"111110101000",
		"011000100001",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001000000000",
		"001100000000",
		"111010011000",
		"111110101001",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110101000",
		"111110010111",
		"101000110001",
		"101000110001",
		"100100110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110010",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"100100100001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"100100110001",
		"100100110001",
		"100100110001",
		"100100110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"101000110001",
		"100100110010",
		"110010011000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110110010111",
		"111110010111",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110010110",
		"111110010110",
		"111110010110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110010110",
		"111110010110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110000110",
		"111110010110",
		"111110010110",
		"111110000110",
		"111101110110",
		"111101010100",
		"111000010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000100010",
		"111100110100",
		"111000110011",
		"111000110011",
		"110101000011",
		"110101000011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111000110011",
		"111001000100",
		"111001000100",
		"111000110010",
		"111000100001",
		"111100110001",
		"111000100010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000100010",
		"111000110010",
		"111000110010",
		"111000100001",
		"111000110010",
		"111000110010",
		"111000100001",
		"111000100001",
		"111100110010",
		"101100000000",
		"101100000001",
		"101000000001",
		"101100000001",
		"101100000000",
		"101100000000",
		"101100000000",
		"101100000000",
		"101100000000",
		"101100000000",
		"101100000000",
		"101100000000",
		"101000000000",
		"101000000001",
		"101100010001",
		"101100010001",
		"101000000000",
		"111000110010",
		"111000110001",
		"111100100001",
		"111000110001",
		"111000110001",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110010",
		"111000110001",
		"111000110010",
		"111000110010",
		"111000110010",
		"110000010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010001",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010001",
		"110100010001",
		"110000010000",
		"110000010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110000010001",
		"101100100001",
		"110110001000",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111011101101",
		"110111001010",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110101000",
		"111101100101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000001",
		"111100000001",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000001",
		"111000000001",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"110000010001",
		"111010000111",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111101100101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111110111000",
		"111110111000",
		"111101110101",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111101100101",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111101100101",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111011001000",
		"111010111000",
		"111110111000",
		"111101110101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111101110101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111101110101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000000",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111101100101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111010001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111101100100",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111001111000",
		"111111101111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110110111010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111110111000",
		"111110101000",
		"111101100101",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001000",
		"111111101111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110110111010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111111001001",
		"111110111000",
		"111110111000",
		"111101110101",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"110101111000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111101100101",
		"110100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110000000000",
		"110110001000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111101110101",
		"111000010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111010001000",
		"111111111110",
		"111111111110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110110111010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111001",
		"111110111000",
		"111001110101",
		"110100010000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000001",
		"111000000001",
		"111000000001",
		"111000000000",
		"111000000000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"111100000001",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"111000000000",
		"110000010001",
		"110101111000",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111110111001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111000",
		"110101110101",
		"110000100001",
		"110100010000",
		"110000010000",
		"110000010000",
		"110000010000",
		"110000010000",
		"110000010000",
		"110000010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110100010000",
		"110000010000",
		"110000010001",
		"110000010000",
		"110000010000",
		"110000010001",
		"110000010001",
		"110000010001",
		"101100010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"101100010001",
		"101100010001",
		"110000010001",
		"101100010001",
		"110000100010",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"101100010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110100010001",
		"110100000000",
		"111000010000",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000000000",
		"110100010000",
		"110100010001",
		"101100010000",
		"101100010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"110000010001",
		"101100010001",
		"101100010010",
		"101100010010",
		"101100100001",
		"101100100001",
		"101100010001",
		"110000010001",
		"110000010001",
		"101100100010",
		"110110001001",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"111011001010",
		"111011001001",
		"111110111000",
		"111110111000",
		"111110111000",
		"111011001001",
		"111011001001",
		"111111001001",
		"111111001000",
		"111110111000",
		"111110111001",
		"111111001001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111110111001",
		"111111001001",
		"111110111001",
		"111110111001",
		"111110111000",
		"111110010111",
		"111110011000",
		"111110010111",
		"111110100111",
		"111110010111",
		"111110010111",
		"111110010111",
		"111110010111",
		"111110010111",
		"111110010111",
		"111110010111",
		"111110011000",
		"111110011000",
		"111110101000",
		"111110011000",
		"111110011000",
		"111110101010",
		"111111001011",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001101",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001011",
		"111110111011",
		"111100110011",
		"111000010001",
		"111100010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100010000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111000000000",
		"111000010001",
		"111101010101",
		"111110111011",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111001100",
		"111111101110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111110111001",
		"111010111010",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101110",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100000001",
		"111101010110",
		"111111101110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101101",
		"110111001010",
		"111010111001",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111001",
		"111010111001",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111001",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111110111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111110111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111000",
		"111010111001",
		"110111001011",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111101111",
		"110100110011",
		"111000000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"111100000000",
		"110100010001",
		"111001100110",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111",
		"111111111111");
	-- Le nombre de vecteur : 60160
	
BEGIN
	PROCESS (RST, HCOUNT, VCOUNT)
	BEGIN
		IF (RST = '1') THEN
			RED <= (OTHERS => '0');
			GREEN <= (OTHERS => '0');
			BLUE <= (OTHERS => '0');
		ELSE
			-- correspondance des pixel
			IF (HCOUNT < XMAX AND VCOUNT < YMAX) THEN
				RED <= data_vector((to_integer(IEEE.NUMERIC_STD.unsigned(VCOUNT)) * XMAX) + (to_integer(IEEE.NUMERIC_STD.unsigned(HCOUNT))))(3 DOWNTO 0);
				GREEN <= data_vector((to_integer(IEEE.NUMERIC_STD.unsigned(VCOUNT)) * XMAX) + (to_integer(IEEE.NUMERIC_STD.unsigned(HCOUNT))))(7 DOWNTO 4);
				BLUE <= data_vector((to_integer(IEEE.NUMERIC_STD.unsigned(VCOUNT)) * XMAX) + (to_integer(IEEE.NUMERIC_STD.unsigned(HCOUNT))))(11 DOWNTO 8);
			ELSE
				RED <= (OTHERS => '0');
				GREEN <= (OTHERS => '0');
				BLUE <= (OTHERS => '0');
			END IF;
		END IF;
	END PROCESS;
END rtl;