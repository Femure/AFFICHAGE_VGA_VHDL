LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY terrain_aff IS
    PORT (
        HCOUNT, VCOUNT : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
        IS_TERRAIN : OUT STD_LOGIC
    );
END terrain_aff;

ARCHITECTURE rtl OF terrain_aff IS
    CONSTANT SCREEN_WIDTH : INTEGER := 640;
    CONSTANT SCREEN_HEIGHT : INTEGER := 480;
BEGIN
    IS_TERRAIN <= '1' WHEN ((HCOUNT > SCREEN_WIDTH/2 - 2 AND HCOUNT < SCREEN_WIDTH/2 + 2) AND VCOUNT <= SCREEN_HEIGHT) ELSE
                '0';
END rtl;