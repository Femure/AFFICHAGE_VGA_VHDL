LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY memory_rom IS
    PORT (
        RST, HCOUNT, VCOUNT, FLAG, XMAX, YMAX : IN STD_LOGIC;
        RED, GREEN, BLUE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        DEP_IMA : OUT STD_LOGIC
    );
END memory_rom;

ARCHITECTURE rtl OF memory_rom IS

    TYPE data_Array IS ARRAY (0 TO 189000) OF std_logic_vector(11 DOWNTO 0);

    -- Initialisation des données
    CONSTANT data_vector : data_Array := (
        "000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000000000",
				"000000010001",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110011",
				"001100110011",
				"001000110011",
				"000100100010",
				"000100100010",
				"000100100010",
				"000000010001",
				"000000000000",
				"000100010001",
				"001000100010",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000100010",
				"001100110011",
				"001101000100",
				"001100110011",
				"001101000100",
				"010001010101",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"001000110011",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"000100100010",
				"000100100010",
				"001101000100",
				"010101100110",
				"010101100110",
				"010001100110",
				"010101100110",
				"010101110111",
				"011001110111",
				"010101100110",
				"001101010101",
				"001101010101",
				"010101100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101000100",
				"001000110011",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000000000",
				"000000010001",
				"000100100010",
				"001000110011",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101110111",
				"010101110111",
				"010001100110",
				"001001000100",
				"000100110011",
				"000100100010",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"000000010001",
				"000100100010",
				"000000100010",
				"000000010001",
				"000000010010",
				"000100100010",
				"000100100011",
				"000100100010",
				"000100100010",
				"000000010001",
				"000100010010",
				"001000110011",
				"001101000100",
				"001101000100",
				"010001010110",
				"011001110111",
				"010101110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010000111",
				"010101110111",
				"010001110111",
				"011110011001",
				"011010011001",
				"011010011000",
				"011010001000",
				"010110001000",
				"010110000111",
				"010101110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101111000",
				"010001100110",
				"010001010110",
				"010001010101",
				"010101100110",
				"001101010101",
				"000100110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100100010",
				"000100100010",
				"001000110011",
				"001101000100",
				"010001100110",
				"011001110111",
				"010001100110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"011001111000",
				"011001110111",
				"010101100110",
				"001101000101",
				"010001010110",
				"011001110111",
				"100010011010",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010001000",
				"011010011001",
				"011010101001",
				"011010011001",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010001000",
				"010110011001",
				"011010011001",
				"010110001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"010001110111",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"010001100110",
				"001101010101",
				"001001000100",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110011",
				"000100100010",
				"000100100010",
				"000100100010",
				"000000010001",
				"001000110011",
				"001101000100",
				"001101000100",
				"001001000100",
				"010001100110",
				"010101110111",
				"010101100110",
				"010001100110",
				"010101100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011010001000",
				"011010011001",
				"011010001000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"011010001001",
				"011110011001",
				"011010001000",
				"010001100110",
				"010001110111",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010101110111",
				"010001110111",
				"010110001000",
				"011010101001",
				"011110101010",
				"010110011001",
				"010010000111",
				"010001110111",
				"010010000111",
				"010110001000",
				"011010101001",
				"011010011001",
				"010010001000",
				"010001110111",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010001110111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001000110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000010000",
				"000000000000",
				"000000010001",
				"001000110010",
				"001000110011",
				"001000110011",
				"000000010001",
				"000000010001",
				"000100100010",
				"001100110100",
				"010101100110",
				"010001010101",
				"001101000100",
				"000100100010",
				"000100010001",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"000100010001",
				"000000000001",
				"000000000000",
				"000000000000",
				"001000100010",
				"001101000100",
				"010001010101",
				"001000110011",
				"001000110011",
				"010001010101",
				"011001110111",
				"011001110111",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001100110",
				"011010000111",
				"011010001000",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110011001",
				"011010011000",
				"010101110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011010001000",
				"010110001000",
				"011010001000",
				"011010011000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011110101010",
				"011110101010",
				"010110001000",
				"010001110111",
				"011010011001",
				"011110101010",
				"011010011001",
				"010110001000",
				"010001100110",
				"010101111000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110011000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110001000",
				"010110011001",
				"010110011000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010101010",
				"011010011001",
				"010001111000",
				"001101100111",
				"010001110111",
				"010010001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"010001100110",
				"001101000100",
				"001000110011",
				"000100010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"010001010101",
				"010101100110",
				"010101110111",
				"010101100110",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101110111",
				"011001110111",
				"011010001000",
				"011001110111",
				"010001010101",
				"001101000100",
				"001101010101",
				"010001010101",
				"010001010101",
				"010101100110",
				"001101010101",
				"000100100010",
				"000000010001",
				"000000010001",
				"000100100010",
				"001100110100",
				"010001010101",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010101110110",
				"011001110111",
				"010101110111",
				"011001110111",
				"011010000111",
				"011110001000",
				"011010001000",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010110000111",
				"011010001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110000111",
				"011010011000",
				"011010011000",
				"010110001000",
				"011010011001",
				"011010011000",
				"011010011001",
				"011010011000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010101001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010110001000",
				"011010101010",
				"011010011001",
				"010110001000",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010110001000",
				"011010011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010001110111",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010101010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"010001100110",
				"001101000100",
				"000100100010",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000100010",
				"001001000100",
				"010001100110",
				"010001100110",
				"001001000100",
				"001101010101",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"010101110111",
				"010101100111",
				"010001100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101110111",
				"001101010101",
				"001101010100",
				"010001010110",
				"010101100110",
				"011010001000",
				"011010001000",
				"010101100111",
				"010001100110",
				"010101100111",
				"011110001000",
				"011110011001",
				"011010001000",
				"010101110111",
				"010001100110",
				"011010001000",
				"011110011001",
				"011110011001",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010110001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010011000",
				"010110011000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"011010011001",
				"011010101010",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110011001",
				"010010001000",
				"010110001001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001000",
				"010001110111",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001001000100",
				"000100100010",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000100010",
				"001101010101",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110000111",
				"010001110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001110111",
				"010001100110",
				"001101010101",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010001110111",
				"010001100110",
				"010001100110",
				"010110000111",
				"010110001000",
				"011010001000",
				"010001100110",
				"001101100101",
				"010101110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011010001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"011010011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"010110001000",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010110001000",
				"011010011000",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110000111",
				"010001110110",
				"010001110111",
				"011010011000",
				"011010011000",
				"010110011000",
				"011010011001",
				"011010011001",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010001110111",
				"010110001000",
				"011010101010",
				"011010011001",
				"010010001000",
				"010010001000",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110011000",
				"010110001000",
				"010001110111",
				"010110001000",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010101010",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010001110111",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101000100",
				"000100100010",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100100011",
				"001101000101",
				"010001100111",
				"011010001001",
				"011010011001",
				"010110001000",
				"010110001001",
				"011010011001",
				"010110001000",
				"010001110111",
				"010110001000",
				"010010000111",
				"010001110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010001100111",
				"010001110111",
				"010110001000",
				"011010001000",
				"010110001000",
				"010001100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"011010011001",
				"010110001000",
				"010001110111",
				"010101110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110000111",
				"010110001000",
				"011010011001",
				"011110101001",
				"011010001000",
				"010110000111",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"010001110111",
				"010001110111",
				"011010001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"011010001000",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110000111",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"011010101010",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"011010101010",
				"010110011000",
				"010010000111",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110011000",
				"010110001000",
				"010010000111",
				"010001111000",
				"010110001000",
				"011010011001",
				"011010011010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001001",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110001001",
				"001101111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"001101110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"001101100110",
				"010001100110",
				"001101000101",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100011",
				"001101000100",
				"001101010101",
				"001101010101",
				"010001100110",
				"010101111000",
				"011010001001",
				"010110001001",
				"010010001000",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010001110111",
				"001101100110",
				"010001110111",
				"011010001001",
				"011010001000",
				"010110001000",
				"011010001000",
				"010001100110",
				"010001110110",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110000111",
				"010001110111",
				"010110000111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011110101010",
				"011010011001",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110011001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011000",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010011001",
				"011010001000",
				"010101110111",
				"010101110111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001110111",
				"011010011001",
				"011110101010",
				"011010011001",
				"010110001000",
				"010001110111",
				"011010011001",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010110011001",
				"010110001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110011001",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"001110001000",
				"010010001000",
				"001110001000",
				"001110000111",
				"010010001000",
				"010010000111",
				"001101110111",
				"001101100110",
				"010001100110",
				"010001100110",
				"001001000100",
				"000000010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000110100",
				"010101110111",
				"011010011001",
				"011110011010",
				"011110011010",
				"011010001000",
				"010001110111",
				"010110001001",
				"011010101010",
				"011010011010",
				"001101111000",
				"001101110111",
				"010010001001",
				"010110011001",
				"010110001000",
				"010110011001",
				"010010001000",
				"010001110111",
				"010110001000",
				"010110001000",
				"010001110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"011010101001",
				"011010101010",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011000",
				"011010011001",
				"010110011000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010001000",
				"010001110111",
				"010110000111",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110101010",
				"011010001000",
				"010101110111",
				"011010001001",
				"011010011001",
				"011110011001",
				"011010011001",
				"010110001000",
				"011010011000",
				"010110001000",
				"010001110111",
				"010001110111",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110110",
				"010001110111",
				"010101110111",
				"010001100110",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011000",
				"011010011000",
				"011010011001",
				"011010011000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010110001000",
				"011010011001",
				"010110011001",
				"010001111000",
				"010010001001",
				"010110011001",
				"011010101011",
				"011010101010",
				"010010001000",
				"010110001001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"001101111000",
				"001101111000",
				"010010001001",
				"010110011001",
				"010010001000",
				"010010001000",
				"001101110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000000000",
				"000000000001",
				"001001000100",
				"010110001000",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010011010",
				"010110001000",
				"011010011001",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110011001",
				"010001111000",
				"010001111000",
				"010110011001",
				"011010101010",
				"011010011001",
				"011010001001",
				"010101111000",
				"010001100110",
				"010101110111",
				"011010011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010001001",
				"010110001000",
				"011010011001",
				"011010011001",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"011010101010",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"011010011001",
				"011010101010",
				"011010101010",
				"011110101010",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010001110111",
				"010110000111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110101010",
				"011010011001",
				"011010011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011010011010",
				"010110001001",
				"010110011001",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011001",
				"011110011001",
				"011110101010",
				"010110101010",
				"010010011001",
				"010110011000",
				"001101110110",
				"010110000111",
				"010110011000",
				"010110011001",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101010",
				"010110011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"001101111000",
				"001101111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010001111000",
				"001101100110",
				"001001010110",
				"001001010101",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110100",
				"010001111000",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110101010",
				"010110011001",
				"010001111000",
				"010010001000",
				"010110001001",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010010001000",
				"001101110111",
				"010010001000",
				"010110001001",
				"010110001000",
				"011010001001",
				"011010001000",
				"010101110111",
				"010110001000",
				"011010001000",
				"010001110111",
				"010001110111",
				"001101100110",
				"010101111000",
				"011010011001",
				"011110011001",
				"010110001000",
				"010001100111",
				"010101111000",
				"010110001000",
				"010110001001",
				"011010011001",
				"010110001001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"010110001001",
				"010110001000",
				"011010011001",
				"011010011010",
				"011010011010",
				"011110101010",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011110101010",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011110101010",
				"011010011010",
				"010110001001",
				"011010011001",
				"011010011001",
				"011110101010",
				"011010011001",
				"010110001000",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001000",
				"010110011001",
				"011110101011",
				"011010101010",
				"011010101010",
				"011110111010",
				"011110101010",
				"011010101010",
				"011110101001",
				"011010101010",
				"011010111011",
				"010110101010",
				"011010101001",
				"010110000111",
				"010110000111",
				"010110001000",
				"010010001000",
				"001101111000",
				"010010001010",
				"010110011010",
				"010110001001",
				"010110001001",
				"011010011001",
				"010110001000",
				"010001111000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"001101111000",
				"001101100111",
				"001101100110",
				"001001000100",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100011",
				"001001000101",
				"010001111000",
				"011010011010",
				"010110101010",
				"010110011010",
				"010110101010",
				"011010101010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"010110011001",
				"010001111000",
				"010001110111",
				"010001110111",
				"010101111000",
				"011010001001",
				"011010001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010001110111",
				"010001100111",
				"001101100110",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010001001",
				"010101111000",
				"010001110111",
				"010001110111",
				"011010001001",
				"011110101010",
				"011110101010",
				"010110001000",
				"001101100110",
				"010010001000",
				"011010101010",
				"011110101010",
				"011010011001",
				"010110011001",
				"010110001000",
				"011010011001",
				"010110001001",
				"011010011001",
				"011110011010",
				"011010011001",
				"011110011010",
				"011010011001",
				"010110001000",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110101010",
				"011110101011",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011001",
				"011110011010",
				"010110001000",
				"010001110111",
				"011010011001",
				"011110101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010111011",
				"011111001100",
				"010110101010",
				"011010101001",
				"011110011001",
				"011110101001",
				"010110001000",
				"010001111000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010110001001",
				"011010011001",
				"010110001000",
				"001101110111",
				"010010001001",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010001111000",
				"001101110111",
				"001101100111",
				"010001100110",
				"001000110100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001101010101",
				"010101110111",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010011010",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010001110111",
				"010001110111",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011010",
				"011010101010",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010011001",
				"010110001000",
				"010001110111",
				"011010001001",
				"011010011001",
				"010110001001",
				"011010011001",
				"011010011001",
				"010010001000",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010011001",
				"011010001001",
				"011110011001",
				"011010011001",
				"010101111000",
				"010001111000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010001111000",
				"010110001000",
				"011010001001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010101110111",
				"010110001000",
				"010110001000",
				"011010011000",
				"011010011001",
				"010110001000",
				"010110000111",
				"010110001000",
				"011010011001",
				"011010101010",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011001",
				"011110101010",
				"011010011001",
				"011010011001",
				"010001111000",
				"010010000111",
				"011010101001",
				"011110101010",
				"011110101010",
				"011110101001",
				"010110011001",
				"010010001000",
				"010110001000",
				"010010011001",
				"010110011001",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010101001",
				"011110011000",
				"011110011000",
				"011110001000",
				"010101111000",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"001101111000",
				"001101100111",
				"010001100111",
				"001101010101",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000001",
				"000000000000",
				"000000000000",
				"001101000100",
				"011010001001",
				"011110101010",
				"011010101011",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110101010",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010010001001",
				"010110011010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010011010",
				"010110011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010101111000",
				"010001100111",
				"010110001000",
				"011110101010",
				"011010001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"011010001000",
				"011010011000",
				"011010011001",
				"011110101001",
				"011010101001",
				"010110011001",
				"010110001000",
				"010110011001",
				"011110101011",
				"011010011010",
				"010110011001",
				"010110001001",
				"011010011010",
				"011110101011",
				"010110011001",
				"010110011001",
				"010110001000",
				"010010000111",
				"011010011001",
				"011110101001",
				"011110101001",
				"011110101010",
				"011010011001",
				"010010000111",
				"001101110111",
				"010010001000",
				"010110011001",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010101010",
				"011110111011",
				"011110011000",
				"010001010100",
				"010001010101",
				"011001110111",
				"011001111000",
				"010101111000",
				"001101111000",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010101010",
				"010110101010",
				"011010101011",
				"010110101010",
				"010010001001",
				"001101111000",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"001101111000",
				"001101100111",
				"010001100111",
				"010001100110",
				"001000110100",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"010101110111",
				"011110101010",
				"011010101010",
				"011010111011",
				"010110111011",
				"010010011010",
				"010110101010",
				"011010101011",
				"010110101011",
				"010110011010",
				"011010101011",
				"011010101011",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110101010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010001100111",
				"011110011001",
				"011110011010",
				"010110001000",
				"010001110111",
				"010001100110",
				"010001110111",
				"010001110111",
				"011010011001",
				"011010001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010101001",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110001001",
				"011010011010",
				"011010101011",
				"010110011001",
				"011010011010",
				"011010011010",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011000",
				"011110101001",
				"011110101001",
				"010110001000",
				"001101110111",
				"010010001000",
				"010110101010",
				"011010111011",
				"010110111011",
				"010110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011110111011",
				"011110101001",
				"010001100101",
				"001000110010",
				"001000100001",
				"001100110011",
				"010001000101",
				"011010001000",
				"010001111000",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110101010",
				"011010101010",
				"010110011010",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"001110001001",
				"010010011010",
				"010110011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"010001111000",
				"001101111000",
				"001101100111",
				"010001110111",
				"001101010101",
				"000000010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001101000101",
				"011010011010",
				"011010101011",
				"010110101010",
				"011010111100",
				"010110111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010010001001",
				"010010011001",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010010001000",
				"010110001001",
				"010010001000",
				"011010011010",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"011110101010",
				"011110101010",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010011001",
				"011110101010",
				"011010011001",
				"010001100110",
				"010001110111",
				"011110011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010101010",
				"011010011001",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011001",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"010110011001",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011010011001",
				"010110001000",
				"011010001000",
				"011010011001",
				"010010000111",
				"001101110111",
				"010110011001",
				"010110101010",
				"011010111011",
				"011010111011",
				"010110111100",
				"011010111100",
				"011010111101",
				"011010101100",
				"100010111011",
				"010101110110",
				"001000100010",
				"001000100001",
				"001000010001",
				"001000010001",
				"000100010010",
				"011001110111",
				"010110001001",
				"010110011001",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"001101110111",
				"010001110111",
				"010001100110",
				"000100110011",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001101010101",
				"010110001001",
				"011110101011",
				"010110101011",
				"010010101010",
				"011011001100",
				"010110101011",
				"010110101011",
				"010110011011",
				"010110011010",
				"010110101011",
				"011010101100",
				"010110101011",
				"010010101010",
				"010010101010",
				"010110101010",
				"010010011001",
				"010110101010",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010010001000",
				"010010001001",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110011001",
				"010001111000",
				"001101100111",
				"011010001001",
				"100010101011",
				"011010011001",
				"010110001000",
				"010001110111",
				"010001110111",
				"011110011010",
				"100010101010",
				"010101111000",
				"010101110111",
				"011010011001",
				"011010001001",
				"011010011001",
				"011010001001",
				"010001110111",
				"010001100111",
				"010110001000",
				"011010011001",
				"011110011010",
				"011010001001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010101010",
				"011110101011",
				"011110101010",
				"011010011001",
				"011010011001",
				"011010001001",
				"010101111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010110011001",
				"011010101010",
				"011010101011",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010110011001",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110001000",
				"001101100110",
				"010001110111",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110011001",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010111100",
				"011011001101",
				"011010111101",
				"011010101011",
				"011110101010",
				"010101100101",
				"000100010000",
				"001000010000",
				"001100100001",
				"001100010010",
				"000100000000",
				"001101000100",
				"011010001000",
				"010110001001",
				"010010011001",
				"010010011010",
				"001110001001",
				"010010001001",
				"010010011010",
				"010110011010",
				"010010011010",
				"010010001001",
				"001110001001",
				"010010001001",
				"010010011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"001101110111",
				"001101100111",
				"010001100111",
				"001001000101",
				"000000010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001001000101",
				"010110001001",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"010110101011",
				"011010111100",
				"011110111100",
				"011010101100",
				"010110011011",
				"011010101100",
				"011010101100",
				"010110111011",
				"010010101010",
				"010110111011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110011010",
				"011010101010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010101011",
				"011010101010",
				"010110011010",
				"011010101011",
				"011010101010",
				"010010001000",
				"010110001001",
				"011110101011",
				"100010101011",
				"011110101010",
				"011010011001",
				"010001100111",
				"010001100111",
				"011010001000",
				"011010011001",
				"010110001000",
				"010101111000",
				"010101110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101111000",
				"010110001000",
				"011110011010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011010011001",
				"010110001000",
				"011010001000",
				"011110011001",
				"011110101010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010101010",
				"011010101011",
				"011110111011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110101010",
				"011010011001",
				"010110001000",
				"010110011001",
				"010010001001",
				"010110011010",
				"011010111100",
				"010110011010",
				"011010101100",
				"011110101011",
				"011010001000",
				"010001000011",
				"001000010001",
				"000100000000",
				"010000110010",
				"001100010001",
				"001000000001",
				"000100010001",
				"010001010101",
				"011010011010",
				"010010011001",
				"001110001001",
				"010110101011",
				"010110101011",
				"010010001001",
				"010110011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"001101110111",
				"001101100111",
				"001101010110",
				"000100110011",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"010001111000",
				"011010101010",
				"011010101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101100",
				"011110111101",
				"011010101100",
				"011010101011",
				"010110011011",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110011010",
				"011110111100",
				"100011011110",
				"100011011101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110001001",
				"010110011001",
				"010010001001",
				"010110011001",
				"011110101011",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011001",
				"011010011010",
				"011110101011",
				"100010111011",
				"011010011001",
				"011010011010",
				"010110001000",
				"010101111000",
				"011010011001",
				"100010101011",
				"011110011001",
				"010101111000",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"011010001001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110001001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010011001",
				"010110001000",
				"011010011001",
				"011010101010",
				"011010101010",
				"010110011001",
				"010010001000",
				"010010001001",
				"010110011010",
				"011110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001001",
				"011010011010",
				"010110011010",
				"011110111100",
				"100010101011",
				"010001010100",
				"001100100001",
				"001100100001",
				"000100000000",
				"010000100010",
				"010000100010",
				"001000010001",
				"000100010000",
				"001000110011",
				"010110001000",
				"010110011001",
				"010010001001",
				"010010011010",
				"010010011010",
				"001110001001",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"001110001001",
				"001110001000",
				"010001111000",
				"010001110111",
				"001101100110",
				"001001000100",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100011",
				"010001110111",
				"010110101010",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101100",
				"010110101100",
				"011010111100",
				"011010101100",
				"011010101100",
				"010110011011",
				"011010111100",
				"010110111100",
				"010110111100",
				"010110101011",
				"011010101011",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011001",
				"010001111000",
				"010010001000",
				"010110011010",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110001000",
				"011010011001",
				"011110101010",
				"011010011010",
				"010110001000",
				"010001111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011011",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"011010011010",
				"011010101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"010101111000",
				"001000100010",
				"001000010000",
				"010000110010",
				"000100000000",
				"001100010000",
				"010100110011",
				"010000100010",
				"000100010000",
				"000100010001",
				"010001010110",
				"010110011001",
				"010110011010",
				"010010011010",
				"001110001010",
				"010010001010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110011011",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010001010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011010",
				"001110001001",
				"001110001001",
				"010010001001",
				"010001111000",
				"001101100111",
				"001101010110",
				"001000110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100011",
				"010001100111",
				"011110111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"100110111100",
				"100110101011",
				"001101100110",
				"010110001000",
				"100111011101",
				"011111001101",
				"011110111100",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010101011",
				"011010101011",
				"010110011010",
				"010010001001",
				"010010001000",
				"010010001001",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010011010",
				"010110001001",
				"010110001001",
				"011010011010",
				"100011001100",
				"011110101011",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110001001",
				"011010001001",
				"010110001001",
				"010101111000",
				"011010011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010011011",
				"010110011010",
				"011010011011",
				"011010101011",
				"010110011010",
				"010110011010",
				"011010101011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011110011010",
				"001101000100",
				"001000100001",
				"001100010000",
				"010100110010",
				"000100000000",
				"000100000000",
				"010100110011",
				"011001000011",
				"001000010001",
				"000100000000",
				"001000110100",
				"010110001001",
				"010110011011",
				"010010001010",
				"001110001010",
				"010010011010",
				"010110101011",
				"010110101011",
				"010110011011",
				"010010011010",
				"010010001001",
				"010010011010",
				"010110011011",
				"010110011010",
				"010010001001",
				"001110001001",
				"010010001001",
				"010010001010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010110011010",
				"010010001001",
				"001110001001",
				"010010011010",
				"010010001000",
				"001101100111",
				"010001100110",
				"001101000101",
				"000100010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000000001",
				"001001000101",
				"011010011001",
				"011110111011",
				"011010111011",
				"010110111011",
				"010110111100",
				"011010111100",
				"011111001101",
				"011010111100",
				"011010111100",
				"010110101100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111011",
				"100110101010",
				"011001100101",
				"000100100001",
				"001101000100",
				"011110101010",
				"100111001101",
				"100011001101",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010101011",
				"010110011010",
				"010010011001",
				"010010011001",
				"011010111011",
				"011110111100",
				"011110111100",
				"011010101011",
				"010110011001",
				"010010001001",
				"010110011001",
				"011110111100",
				"011010101011",
				"011010011010",
				"011010101011",
				"010110011010",
				"010010001000",
				"010010001001",
				"011010011010",
				"011010101011",
				"010110011010",
				"010110001001",
				"011010011010",
				"010110001001",
				"010001111000",
				"010001111000",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010001111000",
				"010110011010",
				"011010101010",
				"010110011010",
				"010110001001",
				"010110001010",
				"010010001001",
				"010010001001",
				"010110011010",
				"011010011011",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110001001",
				"010010001001",
				"010110001001",
				"011010101011",
				"011010011011",
				"010110011011",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110001001",
				"011010001001",
				"011110011010",
				"001101000101",
				"001100100001",
				"010000100001",
				"010000110010",
				"001000010000",
				"000100000000",
				"001100100001",
				"011001010011",
				"001100100001",
				"000100010000",
				"000100100010",
				"010101111000",
				"011010011011",
				"010010011010",
				"010010011010",
				"010010101010",
				"010010011010",
				"010110101011",
				"010110011011",
				"010010011010",
				"010010001010",
				"010010001010",
				"010110011010",
				"010010011010",
				"001110001001",
				"010010001001",
				"010010001010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010110011010",
				"010010001001",
				"001110011001",
				"010010011010",
				"001110001000",
				"001101100111",
				"010001100111",
				"010001010110",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000000001",
				"000000000001",
				"001001010110",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011010111100",
				"010110111100",
				"011010111101",
				"011011001101",
				"010110111101",
				"011010111101",
				"011111001110",
				"010110101100",
				"011010111100",
				"011010101100",
				"100010101011",
				"100001110110",
				"001100010000",
				"010000110010",
				"001100110010",
				"001101010100",
				"100010111011",
				"100111001101",
				"100011011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010010011001",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010011010",
				"011010011010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010010001001",
				"010110011010",
				"010110011010",
				"011010101011",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110001001",
				"010110011001",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010001111000",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"011010011011",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011110101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110101011",
				"010010011011",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010110001001",
				"011010011001",
				"001101000100",
				"001100010001",
				"010000100000",
				"010000100010",
				"001100100001",
				"000000000000",
				"000100010000",
				"010101000011",
				"010000100001",
				"001000010000",
				"000100010001",
				"010101100111",
				"011010011011",
				"010110011010",
				"010010011011",
				"010010011010",
				"001110001001",
				"010010011010",
				"010110011011",
				"010110011010",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001001",
				"010010001010",
				"010110011010",
				"010110011010",
				"010010001010",
				"010010001001",
				"010010011010",
				"010010011010",
				"010010001001",
				"010010011010",
				"010010011010",
				"001110001000",
				"001101100111",
				"010001110111",
				"010001100110",
				"000100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010010",
				"010001110111",
				"011110111100",
				"011010111011",
				"010110111011",
				"011011001100",
				"011010111100",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110111100",
				"011011001101",
				"011011001101",
				"010110111100",
				"010110111100",
				"011011001101",
				"011010111100",
				"011110111100",
				"011110101100",
				"011110001001",
				"011001000010",
				"010000010000",
				"011000110010",
				"010000100001",
				"001000110010",
				"011010001000",
				"100010111100",
				"100011001101",
				"011111001110",
				"011010111101",
				"011011001101",
				"011111001110",
				"011010111101",
				"011010111101",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110101100",
				"011110101011",
				"011110111100",
				"011010101011",
				"011010101011",
				"010110011011",
				"010010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011011",
				"011010101011",
				"011110101100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001010",
				"010110011010",
				"011010101011",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010101010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010110101011",
				"010010101011",
				"001110011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"011010011010",
				"010110011001",
				"011010001001",
				"001101000100",
				"001100010001",
				"010000100000",
				"010100110010",
				"001100110010",
				"000000000000",
				"000000000000",
				"010000110010",
				"010100110010",
				"001000010000",
				"000100000000",
				"010001010111",
				"011010011011",
				"010110011010",
				"010010011011",
				"010010011010",
				"001110011001",
				"010010011010",
				"010110011010",
				"010110011011",
				"010110011010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010110011010",
				"010010011010",
				"010010001001",
				"010010011010",
				"010010011010",
				"010010011001",
				"010010011010",
				"010010011010",
				"001110001000",
				"001101111000",
				"010001110111",
				"010001100110",
				"001000110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000101000101",
				"010110011010",
				"011110111100",
				"010110101011",
				"011010111100",
				"011111001101",
				"011010111100",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101100",
				"011011001101",
				"011011001101",
				"010010111100",
				"010110111101",
				"010110111100",
				"011010111101",
				"011110111101",
				"100010111100",
				"011101110111",
				"010000010000",
				"011000110001",
				"010000100000",
				"010000100001",
				"010001000011",
				"010101100101",
				"100010101010",
				"100111011101",
				"100011001110",
				"011010111101",
				"011110111101",
				"100011001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011011001100",
				"011111001101",
				"011110111100",
				"011010101011",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011011",
				"010110011011",
				"010110011011",
				"010010011010",
				"010010001001",
				"011010011011",
				"011010101011",
				"011010011011",
				"011010101011",
				"011110101100",
				"011110101011",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010110001001",
				"010110001010",
				"010110011010",
				"011010011011",
				"011010101011",
				"010110011011",
				"010110011010",
				"010010011010",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101011",
				"010110011010",
				"010110001001",
				"010110001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"010010011011",
				"010010011010",
				"010010011011",
				"010110101100",
				"010010011011",
				"010010011011",
				"001110011010",
				"010010011010",
				"010110011010",
				"010110001001",
				"011010001001",
				"001101000100",
				"010000100001",
				"010000100000",
				"011001000011",
				"010001000011",
				"000000000000",
				"000100000000",
				"010000110001",
				"011001010011",
				"001100010000",
				"000100000000",
				"010001010110",
				"011010001010",
				"010010001010",
				"010010011011",
				"010010011010",
				"010010101010",
				"011010101100",
				"010110011011",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001001",
				"010010001001",
				"010010001010",
				"010010001010",
				"010010011010",
				"010010011010",
				"010010001001",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010011001",
				"010010001001",
				"010001111000",
				"010001111000",
				"010001100111",
				"001001000100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000100010",
				"000100100010",
				"000100110010",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"000100110010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"001000110011",
				"001000110010",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100010001",
				"000100010001",
				"000100100001",
				"000100100001",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010010",
				"010001111000",
				"100010111100",
				"011110111100",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111100",
				"011110111100",
				"011110111100",
				"010110101011",
				"010110101011",
				"011011001101",
				"010110111100",
				"010110111100",
				"010110111101",
				"011011001110",
				"010110111101",
				"011110111100",
				"100010101010",
				"010101000100",
				"010000010000",
				"011000110010",
				"010100110011",
				"010000110011",
				"010000110010",
				"001100110010",
				"011110011000",
				"100111011101",
				"011111001101",
				"100011001110",
				"100111011110",
				"100111011110",
				"011111001110",
				"011010111101",
				"010110111100",
				"010111001100",
				"011011001101",
				"011111001101",
				"011010111100",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110001010",
				"011110111100",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101100",
				"010110011010",
				"010110001001",
				"011010011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"011010101100",
				"011010101011",
				"011010101100",
				"011010101011",
				"010110011010",
				"010010011010",
				"010110011010",
				"010010001010",
				"010010001010",
				"010110011010",
				"010110001010",
				"011110101011",
				"011010011010",
				"010110001001",
				"010110001010",
				"010110011010",
				"011010011011",
				"011010101011",
				"011110101100",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010001001",
				"010110001001",
				"010110001000",
				"010001111000",
				"011010011010",
				"010110001010",
				"010110011010",
				"011010011011",
				"010110011011",
				"010010011010",
				"010010011010",
				"010110011010",
				"010010011010",
				"011010101011",
				"011110111100",
				"011010101011",
				"011010011011",
				"011010011011",
				"010110011010",
				"010010001010",
				"010110001010",
				"011010011011",
				"010110101100",
				"010110101011",
				"010110101100",
				"010110101100",
				"011010101100",
				"010110011100",
				"010110011100",
				"010010011011",
				"001110011011",
				"010010101011",
				"010010011001",
				"010110011001",
				"011010001000",
				"001100110010",
				"010000100000",
				"010100100000",
				"010100110010",
				"011101100101",
				"000000000000",
				"000000010000",
				"010101000010",
				"011001000010",
				"010000100000",
				"001000010000",
				"010001010101",
				"011010011010",
				"010010011010",
				"001010001010",
				"001110011010",
				"010110101011",
				"010010011011",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010110101011",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010110011010",
				"010010011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101000101",
				"000000010010",
				"000000010001",
				"000000010001",
				"000100100010",
				"000100110011",
				"001000110011",
				"001101000100",
				"001101000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001100110",
				"010101100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001100101",
				"010001010101",
				"001101010101",
				"001101000100",
				"001000110011",
				"000100100010",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000000",
				"000100000000",
				"000000000000",
				"000000000001",
				"000100110100",
				"010110011010",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111101",
				"010110111100",
				"010110111100",
				"011010111100",
				"011110111101",
				"011010111100",
				"010110111100",
				"011010111101",
				"011011001101",
				"011010111101",
				"011011001110",
				"011111001111",
				"011010111101",
				"011110111100",
				"011110001000",
				"001100100001",
				"010000100001",
				"010100110010",
				"001000100010",
				"001100100011",
				"010100110010",
				"010000110001",
				"011001110111",
				"100010111011",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011011001101",
				"010111001101",
				"010111001100",
				"010110111100",
				"011011001101",
				"011110111101",
				"011010111100",
				"011010101100",
				"011010011011",
				"011010101100",
				"011110101100",
				"011110111100",
				"011010011011",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101100",
				"011110111100",
				"011010101011",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110001010",
				"010110001010",
				"010110001010",
				"011010101011",
				"011010101011",
				"010110011011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011011",
				"010010001010",
				"010110011011",
				"011010101100",
				"011010011011",
				"011010101100",
				"011010101011",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110011011",
				"011010101100",
				"011010101100",
				"011010101011",
				"010110011011",
				"010110011010",
				"010110001010",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011010",
				"010110001010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010011011",
				"010110011010",
				"010110001010",
				"010110001011",
				"011010011100",
				"011010101100",
				"010110101100",
				"010010101011",
				"010110101100",
				"011010111101",
				"011010101101",
				"011010011100",
				"010110011100",
				"010010011011",
				"001110011010",
				"001110101010",
				"010010011001",
				"010110011000",
				"011001110111",
				"001100100001",
				"010100100001",
				"010000000000",
				"010000100001",
				"011001010100",
				"000000000000",
				"000000000000",
				"010000110001",
				"010100110001",
				"010000100001",
				"001100100001",
				"010101100110",
				"010110011001",
				"001110011010",
				"001110011011",
				"010010011011",
				"010010011011",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010110011011",
				"010110101011",
				"010010011010",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010010011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001100110",
				"001001000101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010011000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011110101010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011110011001",
				"011010011000",
				"011010001000",
				"011010011000",
				"011010011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010000111",
				"011010000111",
				"011010000111",
				"011010000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"010110111100",
				"010110101100",
				"011010111100",
				"011111001101",
				"011110111101",
				"010110111100",
				"010110111100",
				"011010111101",
				"011010111101",
				"011011001110",
				"011011001110",
				"011011001101",
				"011110111100",
				"011001110110",
				"001000100000",
				"010100110001",
				"010101000010",
				"000000000000",
				"001000100010",
				"010101000011",
				"010000100001",
				"011001100101",
				"100110111011",
				"011110111100",
				"011011001101",
				"011110111101",
				"011110111100",
				"011110111101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011010111101",
				"011110111101",
				"011111001110",
				"011111001101",
				"011010111101",
				"011010101100",
				"011010111100",
				"100010111101",
				"011110111100",
				"011010101011",
				"011010011011",
				"010010001010",
				"010010001001",
				"011010101011",
				"011010111100",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110001010",
				"010010001010",
				"010110001010",
				"010110001010",
				"011010011011",
				"011010101100",
				"010110011011",
				"011010101100",
				"011010111101",
				"011010101100",
				"010110011011",
				"010010001010",
				"010110011011",
				"011010101100",
				"011010101011",
				"010110101011",
				"011010101100",
				"011010101100",
				"010110101100",
				"010110101100",
				"010110101100",
				"010110101100",
				"010010101011",
				"010110101011",
				"010110101011",
				"010110011011",
				"010010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010110101011",
				"010110011010",
				"010110011010",
				"011010101011",
				"010110011011",
				"010010001010",
				"010010011010",
				"010110011011",
				"011010101100",
				"010110101100",
				"010010101011",
				"010010101011",
				"010110101100",
				"011010111100",
				"011010101100",
				"011010101100",
				"010110101100",
				"010010011011",
				"001110101010",
				"001110101010",
				"010010011001",
				"010110001000",
				"011001100101",
				"001100100001",
				"010000010000",
				"001100000000",
				"010000100001",
				"010000110011",
				"000000000000",
				"000000010000",
				"010000110001",
				"001100100000",
				"010000100001",
				"001100100010",
				"010101110111",
				"010110011001",
				"001110001001",
				"010010101011",
				"010010011011",
				"010110011011",
				"010010001010",
				"010010001010",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010110011011",
				"010110011011",
				"010010011010",
				"010110011011",
				"010110101011",
				"010110011010",
				"010010001000",
				"001101110111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010101111000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010011001",
				"011110011001",
				"011110101010",
				"011010101001",
				"011010101001",
				"011010101001",
				"011010101010",
				"011010101010",
				"011010101001",
				"011010101001",
				"011010101001",
				"011010011001",
				"011010101001",
				"011010101001",
				"011010101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010101001",
				"011110101001",
				"011110101001",
				"011110011001",
				"011110101001",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101001",
				"011010011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110000111",
				"011010001000",
				"011010000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"001101000100",
				"001000110011",
				"000100100010",
				"000100100001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"010110001001",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011010111101",
				"010110111100",
				"011010111100",
				"011110111101",
				"011010111101",
				"010110111100",
				"010110111101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"100010111100",
				"010101100101",
				"001100110001",
				"010100110001",
				"011001010011",
				"000000000000",
				"001100110011",
				"011101010100",
				"010000100001",
				"011001010100",
				"100110101010",
				"011110111100",
				"011010111101",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011011001110",
				"011111001110",
				"011010111101",
				"011110111101",
				"011111001110",
				"011111001110",
				"011011001101",
				"011010111100",
				"011010111100",
				"011110111101",
				"011110111101",
				"011110101100",
				"011010011011",
				"010110001010",
				"010110001010",
				"010110011011",
				"011010101100",
				"010110101011",
				"010110011011",
				"011010101011",
				"010110011011",
				"010110011010",
				"010110011011",
				"010110011011",
				"011010011011",
				"010110011011",
				"010010001011",
				"010110011100",
				"010110101100",
				"010110011100",
				"010110011011",
				"010110001011",
				"010110001010",
				"010110001010",
				"010110011011",
				"010110011011",
				"011010101100",
				"011010111101",
				"011010111101",
				"011010101100",
				"011010111100",
				"010110101100",
				"010110101100",
				"010010101011",
				"010010011011",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010110011010",
				"010010011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010010011010",
				"010010001010",
				"010110011011",
				"010110101100",
				"010110101011",
				"010010101011",
				"010010101011",
				"010010111011",
				"010010101011",
				"010110101011",
				"011010101100",
				"011010101100",
				"011010101100",
				"010010011011",
				"001110011010",
				"001110011001",
				"010010001000",
				"010101110110",
				"010101010100",
				"010000100000",
				"001100010000",
				"010000010000",
				"010000100010",
				"001100100010",
				"000000000000",
				"000100010000",
				"001100110010",
				"001100100001",
				"001100100001",
				"001100100010",
				"010110001000",
				"010110011010",
				"001110001001",
				"010010011011",
				"010010011010",
				"010110011011",
				"010010001010",
				"010110011011",
				"010110011011",
				"010010011010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010001010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110011011",
				"010110101011",
				"010110011011",
				"010110011011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010001001",
				"001101111000",
				"001101110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010101001",
				"011010101001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110111010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101001",
				"011010011001",
				"011010101001",
				"011010101001",
				"011010101001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011000",
				"011010011000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010000111",
				"010101110111",
				"010001100110",
				"010001010101",
				"001101010100",
				"001001000100",
				"001001000011",
				"000100100010",
				"000100100010",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001001010101",
				"011010101011",
				"011111001101",
				"010110111100",
				"011010111100",
				"010110111100",
				"010110101100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001110",
				"011111001110",
				"011010111101",
				"010110111101",
				"011010111101",
				"011010111101",
				"011110111011",
				"010001010011",
				"010000110001",
				"010101000001",
				"011001100100",
				"000000000000",
				"001101000100",
				"100001100101",
				"010100110001",
				"010101000011",
				"100010001000",
				"100011001101",
				"011010111101",
				"011010111100",
				"011011001101",
				"011111001100",
				"011010111100",
				"011010111101",
				"011111001111",
				"011110111101",
				"011010111101",
				"011010111101",
				"011111001110",
				"011011001101",
				"010110111101",
				"011010111100",
				"011010111101",
				"011110111101",
				"011110101100",
				"011110101100",
				"011010011100",
				"011010011011",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010101100",
				"011010101011",
				"011010011011",
				"011010011011",
				"010110011011",
				"010010001011",
				"010010001010",
				"010110011011",
				"010110011100",
				"010110011100",
				"011010011100",
				"011010011100",
				"011010011011",
				"011010011011",
				"011010011011",
				"010110001011",
				"011010011100",
				"011110101101",
				"011110101101",
				"011010101101",
				"011010101100",
				"010110101100",
				"011010111101",
				"010110101100",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010110011010",
				"011010101011",
				"011010101010",
				"010110011010",
				"010001111000",
				"001101110111",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010101100",
				"010010011011",
				"010010011010",
				"010110011011",
				"010110101100",
				"010110101100",
				"010110011011",
				"010110101100",
				"010110111100",
				"010110111100",
				"010010101011",
				"010010101011",
				"010110101100",
				"011110101101",
				"011110101101",
				"011010011011",
				"010110011010",
				"010110011001",
				"011010001000",
				"011001110110",
				"010101000011",
				"010000100000",
				"010000010000",
				"001100010000",
				"001100010000",
				"010000110010",
				"000000000000",
				"000100010001",
				"001000100001",
				"001100100010",
				"001100100010",
				"010001000100",
				"011010011001",
				"010110101010",
				"001110011010",
				"010010011010",
				"010010001010",
				"010110011011",
				"010010001010",
				"010010001010",
				"010110011011",
				"010110011011",
				"010110011011",
				"010010001010",
				"010010011010",
				"010010011011",
				"010110011011",
				"010110011011",
				"010010011011",
				"010010011011",
				"010110101011",
				"011010101100",
				"011010101100",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101010",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010111010",
				"011110111010",
				"011110111010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011010111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101001",
				"011010101001",
				"011010011001",
				"011010011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"001101010100",
				"001001000100",
				"001000110011",
				"000100110010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"010001111000",
				"011110111100",
				"011011001100",
				"010110111100",
				"011011001101",
				"010110111100",
				"010110101100",
				"011010111101",
				"011010111100",
				"010110101100",
				"010110101100",
				"011010111101",
				"011010111101",
				"011011001110",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011111001101",
				"011110111011",
				"010001000011",
				"010000110001",
				"010100110001",
				"011001010011",
				"000000000000",
				"001100110011",
				"100001110110",
				"011001000011",
				"010100110010",
				"011001100110",
				"100010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011010111100",
				"011110111110",
				"011111001111",
				"011111001110",
				"011010111110",
				"011010111110",
				"011011001110",
				"011010111101",
				"010110111101",
				"010110101100",
				"011010101100",
				"011010111101",
				"011010111101",
				"011010101100",
				"011010101100",
				"011010011011",
				"010110011011",
				"010110011011",
				"011010101100",
				"011010101011",
				"011010101100",
				"011110111100",
				"011010101100",
				"011010101100",
				"011010101100",
				"010110011011",
				"010110011011",
				"010110011011",
				"011010101100",
				"011110101101",
				"011010101100",
				"011010011100",
				"011010011011",
				"011010001011",
				"011010001011",
				"011010001011",
				"011010001011",
				"011110011100",
				"100010101101",
				"100010101101",
				"011110101101",
				"011110101101",
				"011110101101",
				"011110101101",
				"011010101100",
				"010110011011",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010010001010",
				"010010011011",
				"011010111100",
				"011010111101",
				"010110101100",
				"011010101100",
				"011010101100",
				"010110111100",
				"010010111100",
				"010010101011",
				"010010101011",
				"011010101100",
				"011110101101",
				"011110101101",
				"011110101100",
				"011110101100",
				"011110101011",
				"100010011010",
				"011101110111",
				"010100110010",
				"010000010000",
				"001100010000",
				"001100010000",
				"001000000000",
				"010000110010",
				"000100000000",
				"001100100010",
				"001000010001",
				"000100010001",
				"001000100011",
				"010101100111",
				"011010011010",
				"010010011010",
				"001110011010",
				"010010101011",
				"010110011011",
				"010110011010",
				"010110001010",
				"010010001010",
				"010110011011",
				"010110011011",
				"010110011011",
				"010010011011",
				"010010011011",
				"010010011011",
				"010110101011",
				"010110101011",
				"010110011011",
				"010110011011",
				"010110101011",
				"010110101100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111010",
				"011110111011",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111011",
				"011010111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110011000",
				"011010011001",
				"011010011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"010110001000",
				"010110000111",
				"010101110111",
				"010001110110",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001010101",
				"001101000100",
				"001101000100",
				"001000110010",
				"000100100001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"010110001001",
				"011111001100",
				"010110111100",
				"010110111100",
				"011011001101",
				"010110111100",
				"011010111100",
				"011111001101",
				"011011001101",
				"010110111100",
				"011010111101",
				"011010111101",
				"010110111101",
				"010110111101",
				"011010111101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011110111011",
				"010001010100",
				"010000110001",
				"010000100000",
				"010101000010",
				"000000000000",
				"001000100010",
				"100001110110",
				"011101010011",
				"011000110010",
				"010101000100",
				"100010101011",
				"011010111101",
				"011011001101",
				"011011001101",
				"011111001100",
				"011111001101",
				"011111001110",
				"011111001111",
				"011111011111",
				"011111001110",
				"011011001110",
				"011011001110",
				"011010111101",
				"011010111101",
				"010110101100",
				"010110101100",
				"010110111101",
				"011010111101",
				"011010111101",
				"011010101100",
				"010110101100",
				"010110011011",
				"010110001011",
				"010110001010",
				"010010001010",
				"010110011011",
				"011010111100",
				"011010101100",
				"011010101100",
				"011110101100",
				"011010101100",
				"011010011100",
				"011010011100",
				"011110101101",
				"011110101101",
				"011010011011",
				"010110001011",
				"010110001010",
				"010101111010",
				"010101111010",
				"011001111010",
				"100010001100",
				"100110101101",
				"100110101110",
				"100110111110",
				"100010101101",
				"100010011100",
				"100010101101",
				"011110011100",
				"011010011011",
				"011010011011",
				"011010011011",
				"011010011011",
				"011010011010",
				"011010001010",
				"010110001010",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110111011",
				"011010101011",
				"010110011010",
				"011010101011",
				"011010111100",
				"010110101100",
				"010010011011",
				"010110101100",
				"010110101100",
				"011010111101",
				"011010111100",
				"010110101100",
				"010110101101",
				"010110101101",
				"010010101100",
				"010010101100",
				"010010101100",
				"010010101100",
				"010110101100",
				"011010101101",
				"011010011100",
				"011010011100",
				"011010011011",
				"011010011011",
				"011110011010",
				"011001110111",
				"001100100001",
				"001000010000",
				"001100010000",
				"001100010000",
				"001100010000",
				"010000100001",
				"001000010000",
				"010000110011",
				"001000010001",
				"000000000000",
				"001100110100",
				"011010001001",
				"010110011010",
				"010010011010",
				"010010101011",
				"010110101011",
				"011010011011",
				"011010011010",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110101011",
				"010110011011",
				"010010011011",
				"010110101011",
				"010110101100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101100",
				"011010111100",
				"011010111100",
				"011110111100",
				"100011001100",
				"011010111011",
				"010110101010",
				"011010101011",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011111001011",
				"011111001011",
				"011111001011",
				"011110111011",
				"011110111011",
				"011010101010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011110111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010101001",
				"011010101010",
				"011010101010",
				"011010101001",
				"011010011001",
				"011010011001",
				"011010101001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110110",
				"010001100110",
				"001101010101",
				"001000110011",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"010110011010",
				"011111001101",
				"010110111100",
				"010111001101",
				"011011001101",
				"010110111100",
				"011010111100",
				"011111001101",
				"011011001101",
				"011010111100",
				"011011001110",
				"011111001110",
				"011011001110",
				"010110111101",
				"010110111100",
				"011111001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011110111011",
				"010101100100",
				"010000110001",
				"010000100000",
				"011001000010",
				"000100010001",
				"000100010001",
				"100001100101",
				"011101010011",
				"011000110010",
				"010100110011",
				"011110011010",
				"011010101100",
				"011010111101",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001111",
				"011011001111",
				"011111011111",
				"011011001111",
				"011011001110",
				"011011001110",
				"011010111110",
				"011010111101",
				"011010111101",
				"011010111101",
				"010110101100",
				"011011001110",
				"011111001110",
				"011010111101",
				"011010111101",
				"011010101100",
				"010110011011",
				"010110001010",
				"010010001001",
				"010010011010",
				"011110111100",
				"011010101100",
				"011110101100",
				"011110111101",
				"011010101100",
				"011010011011",
				"011010101100",
				"011110111101",
				"011110101100",
				"011010011011",
				"011010011011",
				"011110011100",
				"011110011011",
				"011110001011",
				"011101111010",
				"100110101101",
				"101110111110",
				"101111001111",
				"101010111110",
				"100010101101",
				"011110001011",
				"011110011011",
				"011010001011",
				"011010001011",
				"010110001010",
				"010110001010",
				"010110001001",
				"010110001001",
				"010110001010",
				"010110001010",
				"010110011010",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"010110011010",
				"010010001001",
				"011010101011",
				"011010101100",
				"010110011011",
				"010110101100",
				"011010111110",
				"011111001110",
				"010110101100",
				"010110101100",
				"011010111101",
				"010110101100",
				"010110101100",
				"010010011100",
				"010010011100",
				"010110101100",
				"011010101101",
				"011010101100",
				"010110011100",
				"010110011100",
				"010110011011",
				"010110011011",
				"010110011010",
				"011110011010",
				"010101110111",
				"001000100010",
				"001000010000",
				"001100010000",
				"001100010000",
				"010000010000",
				"010100100010",
				"001100010001",
				"001100010001",
				"000100000000",
				"000100010010",
				"010001010110",
				"011110011010",
				"010110011010",
				"010010101011",
				"010110111100",
				"010110101011",
				"011010011011",
				"011010011011",
				"011010011011",
				"011010101100",
				"011010101100",
				"010110101100",
				"010110101100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101100",
				"010110101100",
				"010110101100",
				"010110101100",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111011",
				"100011001100",
				"011110111011",
				"011010101010",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011010111010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110000111",
				"011001110111",
				"010101110111",
				"010101100110",
				"010001100101",
				"001101000100",
				"001000110011",
				"000100100010",
				"000000010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000010001",
				"000000010000",
				"000000010001",
				"000100100001",
				"001000100010",
				"001000110010",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"001101000011",
				"001001000011",
				"001000110011",
				"001000110011",
				"001100110011",
				"001101000100",
				"001101000100",
				"010001000101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001100101",
				"010001010101",
				"001101010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"001101000100",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"000100100010",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000010001",
				"000000010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000100011",
				"010110011001",
				"011111001101",
				"011010111100",
				"010111001100",
				"011011001101",
				"011010111100",
				"011010111101",
				"011010111100",
				"011011001101",
				"011010111101",
				"011010111110",
				"010110111101",
				"011011001110",
				"011011001110",
				"011010111100",
				"010110101100",
				"011110111101",
				"011110111101",
				"011010111100",
				"011110111011",
				"011001110110",
				"001100100001",
				"010100100001",
				"100001010100",
				"001000010001",
				"000000000000",
				"011001010100",
				"011001000010",
				"011101010011",
				"010100110011",
				"010101100111",
				"011110101100",
				"011111001101",
				"011010111101",
				"100011011101",
				"011111001101",
				"011011001110",
				"010111001111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011011001110",
				"011010111101",
				"011010111110",
				"011010111110",
				"011010111101",
				"010010101100",
				"010110111101",
				"011111011111",
				"011111011111",
				"011111001110",
				"011010111101",
				"011010101100",
				"010110011011",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110011011",
				"010110011010",
				"010110011010",
				"011010011011",
				"011010101100",
				"011010101100",
				"011010101011",
				"011110101100",
				"011110111101",
				"011110101100",
				"100010101100",
				"100010101100",
				"100010101100",
				"011110011011",
				"100110101101",
				"100110111101",
				"100110101101",
				"100010101100",
				"011110011100",
				"011010011011",
				"011010011011",
				"011010011011",
				"011010011011",
				"010110011011",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010111011",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101100",
				"010110101100",
				"010110101101",
				"011010111101",
				"011010111101",
				"010110101100",
				"010110101011",
				"010110101100",
				"010010101100",
				"010010101100",
				"010110101100",
				"011010101011",
				"011110101100",
				"011110101100",
				"011110011100",
				"011010011011",
				"010110011011",
				"001110011010",
				"010010101011",
				"010010101010",
				"010110011001",
				"011010001000",
				"001100110011",
				"001100100001",
				"001100010000",
				"001100010000",
				"001100000000",
				"010000010000",
				"001100010000",
				"001000000000",
				"000100010001",
				"001000110011",
				"011110011010",
				"011110101011",
				"011010101011",
				"010110111100",
				"011011001101",
				"011010111100",
				"011010011011",
				"011110101011",
				"011010101100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"010110101100",
				"010110111100",
				"011010111101",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"100011001100",
				"100010111100",
				"011110111011",
				"011110111011",
				"100011001100",
				"011110111100",
				"011010101011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110111011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011000",
				"011010001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001010101",
				"001101000100",
				"001100110011",
				"001000110011",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"000100010010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"001000100010",
				"001000100010",
				"001000110011",
				"001000110011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010101",
				"010001010101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011010001000",
				"011010001000",
				"011001110111",
				"011010000111",
				"011010000111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"010101110110",
				"010101100110",
				"010101110110",
				"010101110110",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010001100110",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000100",
				"001101000100",
				"001000110011",
				"001000100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000000001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"010010001001",
				"011111001101",
				"011011001100",
				"010111001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011111001110",
				"011011001110",
				"011011001110",
				"010110111101",
				"011010111100",
				"011110111101",
				"011111001110",
				"011110111101",
				"011010111100",
				"011110111100",
				"011110011000",
				"010000110010",
				"010000010000",
				"010100110010",
				"010101000011",
				"000000000000",
				"010101000011",
				"011101010011",
				"011101000011",
				"011001000011",
				"011001100111",
				"100010101011",
				"011110111101",
				"011110111100",
				"100011001101",
				"100011011110",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111001110",
				"011111001110",
				"011111001110",
				"011011001110",
				"010110111101",
				"011010111101",
				"011010111101",
				"011011001110",
				"011111001110",
				"011110111101",
				"011010111101",
				"011110111101",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110011011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"100010101100",
				"100010101100",
				"011110011011",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011010101100",
				"011010101100",
				"010110011011",
				"010110101011",
				"010110011011",
				"010110011010",
				"010110101010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110101010",
				"011010111011",
				"011010101010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110101100",
				"010110101100",
				"010110101100",
				"010110101100",
				"010110011011",
				"010110011011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010011010",
				"011010011010",
				"011001111001",
				"011001101000",
				"011001111001",
				"011110011010",
				"011010101011",
				"010010011010",
				"010010101010",
				"010010101010",
				"010010011001",
				"011010011001",
				"010001000100",
				"001000010000",
				"001100100001",
				"010000110001",
				"010000100001",
				"010000100000",
				"001000000000",
				"001000010001",
				"001100110011",
				"010001010101",
				"011110011010",
				"011110101011",
				"011010101100",
				"010110111100",
				"011011001101",
				"011010111100",
				"011110101100",
				"011110101100",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111101",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011110111100",
				"100111001100",
				"100111001100",
				"100010111100",
				"100010111100",
				"100011001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011110101011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001110111",
				"010101110111",
				"010101100110",
				"010001010101",
				"001101000100",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001000100010",
				"001000100011",
				"001100110100",
				"010001000101",
				"010001010101",
				"010101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110111",
				"011001110111",
				"011110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101111000",
				"010101111000",
				"011001111000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"011110011000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010000111",
				"011001110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001100110011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000010000",
				"000000010000",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000100011",
				"010110011010",
				"011111001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011010111101",
				"011111001110",
				"011010111110",
				"011011001110",
				"011011001101",
				"011111001101",
				"100011001110",
				"011110111101",
				"011010111101",
				"011010111101",
				"011111001101",
				"100010101010",
				"010001000011",
				"010000100001",
				"010000010001",
				"011101010100",
				"001000010000",
				"001100100001",
				"011101100101",
				"011101000011",
				"011001010011",
				"011001010110",
				"100010011010",
				"100010111100",
				"100010111101",
				"100011001101",
				"100011011110",
				"011111011111",
				"011111101111",
				"011111011111",
				"100011011110",
				"100011011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"011010111101",
				"011010101101",
				"100011011111",
				"100011011111",
				"011010111101",
				"011011001101",
				"011011001100",
				"011010111100",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010011011",
				"011110101011",
				"011110101100",
				"011010011011",
				"011010011011",
				"011010011010",
				"011010011011",
				"011010101100",
				"011010101100",
				"011010101011",
				"011010101100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010010011001",
				"001110001000",
				"001110001000",
				"010010011001",
				"010110101010",
				"011010111011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010010011011",
				"010110101100",
				"010110101100",
				"010010011100",
				"010010011011",
				"010110011011",
				"010110011011",
				"011010011010",
				"100010101011",
				"011010001000",
				"010101100110",
				"010101010101",
				"010101000101",
				"010100110100",
				"010101000101",
				"011101111000",
				"011010001000",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110011001",
				"011110101010",
				"010101100110",
				"000100010001",
				"001000100001",
				"001100110010",
				"010000100001",
				"010000100001",
				"001000010000",
				"001100110010",
				"010101010101",
				"011010001000",
				"100010101011",
				"100010111100",
				"011110111101",
				"011011001101",
				"011111011101",
				"011111001101",
				"100010111101",
				"100010111101",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010111101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011110111100",
				"011110111100",
				"011111001100",
				"100011001100",
				"100011001100",
				"101011011101",
				"101011011101",
				"100111001100",
				"100111001100",
				"100111001101",
				"100011001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011001",
				"011010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101100110",
				"001101010101",
				"000100110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000010010",
				"000100100010",
				"001000110011",
				"001101000101",
				"010001010101",
				"010101100110",
				"010101100110",
				"011001110111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011010001000",
				"011001110111",
				"010101110111",
				"011001110111",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011010011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000100010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000101000101",
				"011010111011",
				"011111011101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011111001110",
				"011111001110",
				"011011001101",
				"011010111110",
				"011010111110",
				"011011001110",
				"011111001110",
				"011010111100",
				"011111001101",
				"011110111101",
				"011010111101",
				"010110111101",
				"011111001101",
				"011110101011",
				"010101100110",
				"001100100010",
				"010000100001",
				"011001000010",
				"011001000010",
				"001100010000",
				"011001010011",
				"011101010011",
				"011001000011",
				"010101000100",
				"011101111000",
				"100110111100",
				"100111001101",
				"100111001101",
				"100011001110",
				"011111001110",
				"011111001111",
				"100011011111",
				"100011001110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111101",
				"011111001110",
				"100011011111",
				"100111011111",
				"101011101111",
				"100111011111",
				"011110111101",
				"011111001110",
				"100011011111",
				"011111001110",
				"011111011110",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010101011",
				"010110011011",
				"010110011011",
				"011010101011",
				"011010101100",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010011011",
				"011010011011",
				"010110011010",
				"011010011011",
				"011010101100",
				"011010101100",
				"010110101011",
				"010110101011",
				"010010101011",
				"010110101011",
				"010010101010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010010011010",
				"010110101011",
				"011010111011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101100",
				"010110101100",
				"010110101100",
				"010110011100",
				"010110011011",
				"011010011011",
				"011110011011",
				"011110011010",
				"100010001001",
				"010101010101",
				"010000100010",
				"010000110010",
				"010100110010",
				"010100110010",
				"011000110011",
				"011001010101",
				"011001100110",
				"011110001000",
				"011110011001",
				"011110101010",
				"011110011001",
				"100010101010",
				"100010011010",
				"010001100110",
				"001000110011",
				"001000100010",
				"001000010000",
				"001000100000",
				"001000010000",
				"001100110010",
				"010101100110",
				"011110011010",
				"100110111101",
				"100010111101",
				"100011001101",
				"011111001101",
				"011111011110",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011011101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011011001101",
				"011111001101",
				"011011001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"100011001100",
				"100011001101",
				"100111011101",
				"100111011101",
				"101111011101",
				"101111011101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"001101010101",
				"000100110011",
				"000000010010",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"000100100010",
				"001000110011",
				"001000110011",
				"001001000100",
				"001101000101",
				"001101010101",
				"010001100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011110011001",
				"011110011001",
				"100010101011",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010011000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"011010000111",
				"011010000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001000100",
				"001101000100",
				"001101000011",
				"001000110011",
				"001000100010",
				"000100100010",
				"001000100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001010110",
				"011111001100",
				"011111001101",
				"010111001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001110",
				"011011001110",
				"011111001110",
				"011011001110",
				"011010111101",
				"010110101011",
				"011010101011",
				"011110111101",
				"011010111101",
				"010110111101",
				"011011001101",
				"011110111100",
				"100010101010",
				"001101000011",
				"001100100001",
				"010100110001",
				"011101010011",
				"010000100001",
				"010000100001",
				"011001000011",
				"011001000011",
				"010000110010",
				"011001010101",
				"100010101011",
				"100110111101",
				"100010111101",
				"100010111101",
				"011110111101",
				"011110111110",
				"100111011111",
				"100111001110",
				"100011001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010101100",
				"011110111101",
				"100011001110",
				"100011001110",
				"100011001110",
				"011110111101",
				"011111001110",
				"100011011111",
				"100011101111",
				"011111011110",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011010101100",
				"011010101011",
				"010110101011",
				"011010101100",
				"011010101100",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010101011",
				"011010011011",
				"011010011011",
				"011010101100",
				"011010111100",
				"011010101100",
				"010110101011",
				"010110101100",
				"010110011011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111100",
				"011010111101",
				"010110101100",
				"010110011100",
				"010110011100",
				"010110011011",
				"011010011011",
				"100010101011",
				"100110011010",
				"011001000101",
				"011000110011",
				"010100100010",
				"011000110010",
				"011000110010",
				"011000110001",
				"011000110010",
				"011101010100",
				"100101100110",
				"101010001001",
				"100110001001",
				"100110011010",
				"100010011010",
				"100010111011",
				"100111001101",
				"100010111011",
				"011010011010",
				"010101111000",
				"010001010101",
				"010101010101",
				"010001010100",
				"011001110110",
				"011110011001",
				"100110111100",
				"100110111101",
				"100010111101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"100010111100",
				"100111001100",
				"101011011101",
				"101011011101",
				"101011011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"100111001100",
				"100011001100",
				"100011001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"001101010101",
				"001001000100",
				"000100110011",
				"000000010010",
				"000000010001",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000010001",
				"000100100010",
				"001000110010",
				"001101000100",
				"010001010101",
				"010101100110",
				"011001110111",
				"011001110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110101010",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010110001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"001000100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000100000001",
				"000000000001",
				"000000010010",
				"001101100111",
				"011111001100",
				"011011001101",
				"010111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011010111110",
				"011111001110",
				"011011001110",
				"011010111101",
				"011110111100",
				"011010101011",
				"011010101100",
				"010110111101",
				"010111001110",
				"011011011111",
				"011110111101",
				"100111001100",
				"010101110111",
				"001000100001",
				"010100110001",
				"011000110001",
				"011001000011",
				"010000100010",
				"010101000010",
				"010100110010",
				"010101000010",
				"010101010100",
				"100010011010",
				"100010101100",
				"100010101100",
				"100010111101",
				"011110101101",
				"011110111101",
				"100111001110",
				"100010111101",
				"100010111101",
				"100010111101",
				"100010111101",
				"011110101100",
				"011110101100",
				"011110101100",
				"100010111101",
				"011110101100",
				"011110101101",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111011111",
				"011111001110",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011010111100",
				"011010101100",
				"011010101100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010011011",
				"010110011011",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010101100",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011110111100",
				"010110101011",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011111001101",
				"011010111101",
				"010010011011",
				"010010011011",
				"010110011100",
				"011010011011",
				"011110011011",
				"100010011011",
				"100010001001",
				"011100110100",
				"011100110011",
				"011100110010",
				"011000110001",
				"011000110001",
				"011000110001",
				"011001000010",
				"011101000011",
				"100101100110",
				"101110001001",
				"101010001001",
				"101010011011",
				"100110101011",
				"100010111100",
				"100011001101",
				"011111001101",
				"100011001110",
				"100111001110",
				"100110111011",
				"100110111010",
				"100110111010",
				"101011011100",
				"100111001101",
				"100111001101",
				"100111001110",
				"100010111101",
				"100011001101",
				"100011001101",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"100011001100",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001100",
				"100111001100",
				"100111001100",
				"101011011101",
				"101111011101",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100011001100",
				"100011001100",
				"011110111100",
				"010110101011",
				"010110101011",
				"010110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001110111",
				"010001110111",
				"001101010110",
				"001001000100",
				"000100110011",
				"000100100010",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101100110",
				"010101100110",
				"010101110110",
				"011001110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011110111010",
				"011110111010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010101010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010110001000",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001000100",
				"001101000100",
				"001101000100",
				"010001000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"001000100011",
				"001000100011",
				"000100110011",
				"010110001001",
				"011111001100",
				"011011011101",
				"011011011101",
				"010111001101",
				"011011001101",
				"011111001110",
				"011111001110",
				"100011011111",
				"011111011110",
				"011111011110",
				"011011001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"100011001101",
				"011110111100",
				"011010101100",
				"011010111110",
				"011011011111",
				"011011011111",
				"011111001101",
				"100011001101",
				"100011001011",
				"010001100101",
				"011001000001",
				"010100100000",
				"011001000010",
				"011000110011",
				"010100110010",
				"010101000010",
				"010101000010",
				"010101000011",
				"100010001001",
				"100110101100",
				"100010101100",
				"100010101101",
				"100010101100",
				"011110101100",
				"011110101100",
				"011010011011",
				"011010011010",
				"011010011011",
				"011110011011",
				"100010101100",
				"100010101100",
				"011110101100",
				"011110011100",
				"011110111101",
				"100011001110",
				"100011011111",
				"011111001110",
				"011010111101",
				"011010111101",
				"100011011111",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100111011111",
				"100011011110",
				"100011001110",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101100",
				"010110101011",
				"010110101011",
				"010110011011",
				"010110011011",
				"011010101100",
				"010110101100",
				"010110101100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"100011001100",
				"100011001100",
				"011110111100",
				"011110111100",
				"011110111101",
				"010110101100",
				"010010011011",
				"010010011011",
				"010110011100",
				"011010011011",
				"011110011011",
				"100010011010",
				"011101100111",
				"100001100110",
				"100001010100",
				"011101000011",
				"011000110001",
				"011000110001",
				"011001000001",
				"011001000001",
				"011001000010",
				"011101010101",
				"101010001001",
				"101010011010",
				"101010101100",
				"100110111101",
				"100010111101",
				"010110111101",
				"010111001101",
				"011010111110",
				"100011001110",
				"100011001101",
				"100111001100",
				"100111001100",
				"100111011100",
				"100011001100",
				"011110111100",
				"100111001110",
				"100010111110",
				"100111001101",
				"100011001101",
				"100011001100",
				"100011001101",
				"100111011101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100111011110",
				"100111011101",
				"100111011101",
				"101011001101",
				"101011001101",
				"101011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100011001100",
				"100011001101",
				"011110111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001010110",
				"001101000101",
				"001000110011",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110011",
				"001101000100",
				"010001010101",
				"011001110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010011001",
				"011110011001",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101010",
				"011110101011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010101111000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001000100",
				"010001000100",
				"010001010100",
				"010001010101",
				"010101010101",
				"010101010101",
				"010001010101",
				"010001010101",
				"001101010110",
				"011110101011",
				"011111001101",
				"100011101110",
				"011111101110",
				"010111001101",
				"011011001101",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011111",
				"100011011111",
				"100011011111",
				"011111001110",
				"010110101100",
				"011010101011",
				"011110111101",
				"011110111101",
				"100011011111",
				"011111011111",
				"010110111101",
				"011111001101",
				"100011001101",
				"101011101110",
				"100111001010",
				"011001100100",
				"011000110001",
				"010000100001",
				"010100110010",
				"010101000011",
				"011101010100",
				"010000110010",
				"010000110011",
				"011110001001",
				"100110111100",
				"100110101100",
				"100110111101",
				"100010101011",
				"100010011011",
				"011010001001",
				"010101111000",
				"010101100110",
				"010101010110",
				"011001101000",
				"100010001001",
				"100010011011",
				"100010101011",
				"100010101100",
				"100010111110",
				"011110111101",
				"011110111110",
				"100011011111",
				"100011011111",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011010111101",
				"010110101100",
				"010110101011",
				"010110011011",
				"010110011011",
				"010110101100",
				"010110101100",
				"010110101100",
				"011010111101",
				"011011001101",
				"011010111101",
				"010110111101",
				"011010111101",
				"011010111101",
				"010110101100",
				"010010101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011010101011",
				"011010101100",
				"010110011100",
				"010010011011",
				"010110011100",
				"010110011100",
				"011010011011",
				"100010101100",
				"100010011010",
				"011001100111",
				"100001100110",
				"100101010101",
				"100001010100",
				"100001010011",
				"011101000010",
				"011001000010",
				"011001000010",
				"011001000011",
				"011001010101",
				"101010011001",
				"101010101011",
				"100110101100",
				"011110111101",
				"011111001110",
				"011011001101",
				"011111011111",
				"011111011111",
				"011111001111",
				"100011001101",
				"100011011101",
				"100011001100",
				"100011001100",
				"100011001100",
				"100111011110",
				"100111001110",
				"100010111101",
				"100111001101",
				"100111001101",
				"100011001100",
				"100011011100",
				"100111011101",
				"100111001100",
				"100111011101",
				"100111001100",
				"100011001100",
				"100111001101",
				"100111011101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011101",
				"101011011110",
				"101111011110",
				"101011011101",
				"101011001100",
				"101011001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100011001100",
				"100011001101",
				"011111001100",
				"010010101010",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101010",
				"010010011001",
				"010010011010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110001000",
				"011010001001",
				"010110001000",
				"010101110111",
				"010101100111",
				"010001100110",
				"001000110100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000010001",
				"000100100010",
				"000100110011",
				"001001000100",
				"001001010101",
				"010001100110",
				"010001110111",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"011010011010",
				"011110101011",
				"100010111100",
				"100010111100",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010001110111",
				"001101010110",
				"001101100110",
				"010101100111",
				"011010001000",
				"011110001001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110110",
				"010001110111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001010110",
				"010001100110",
				"010101100110",
				"010101100111",
				"011001100111",
				"010101100110",
				"010101100110",
				"010101010110",
				"010101010110",
				"010101010101",
				"010101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101100110",
				"010001100111",
				"100010111100",
				"011111001101",
				"100111101111",
				"100011011110",
				"011011001101",
				"011111011110",
				"011111011110",
				"011111001110",
				"100011011111",
				"011111011110",
				"100011011111",
				"100111111111",
				"100111101111",
				"011111011110",
				"011011001101",
				"011010111100",
				"011010111101",
				"011111001101",
				"100011011110",
				"100011011110",
				"011111001101",
				"100011001101",
				"100111011101",
				"101011101110",
				"101011011101",
				"100110101010",
				"011001100110",
				"010001000011",
				"010000110011",
				"010101000100",
				"010000110100",
				"010101000101",
				"100010001001",
				"110011011110",
				"100110111100",
				"100110111100",
				"101011001100",
				"100110111011",
				"100010011001",
				"100010000111",
				"011101100101",
				"100001010101",
				"100001010101",
				"100001010101",
				"011101010101",
				"011101100111",
				"100010001001",
				"100110101100",
				"100110111101",
				"011110111101",
				"011010111101",
				"011111001110",
				"011111011111",
				"100011011111",
				"100111011111",
				"100111011111",
				"101011011111",
				"101011101111",
				"100111011111",
				"100010111101",
				"011110111101",
				"100011001101",
				"100011001110",
				"011011001101",
				"011011011110",
				"011011001101",
				"011111011110",
				"011111001101",
				"010110101011",
				"010110101100",
				"010110101100",
				"010110111100",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111100",
				"010110101100",
				"010110101100",
				"010110111100",
				"010110101100",
				"010010011011",
				"010010011011",
				"010110111100",
				"011010111101",
				"011111001101",
				"011111001110",
				"011011001101",
				"011010111101",
				"011010111101",
				"100011001110",
				"100111001101",
				"100010101100",
				"011110101011",
				"011010011011",
				"010110001011",
				"010110011100",
				"010010011100",
				"010110011101",
				"010110011100",
				"011010011100",
				"100010101100",
				"100010011011",
				"011001100111",
				"011101010101",
				"101001110110",
				"100101010100",
				"011101000010",
				"100001000010",
				"011101000010",
				"011000110001",
				"011001010100",
				"100010001000",
				"100110101011",
				"101011001101",
				"100010111101",
				"011110111101",
				"011110111101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011101",
				"011111011101",
				"011111001100",
				"011111001100",
				"100011011100",
				"100111011101",
				"100111011101",
				"101011011110",
				"101011011110",
				"101011001101",
				"100111001100",
				"100111001100",
				"101011011101",
				"101011011101",
				"100111001100",
				"101011001100",
				"100110111100",
				"101011001100",
				"101011011101",
				"101011001101",
				"100111001100",
				"101011001100",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111011101",
				"100111001101",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101010",
				"010010011010",
				"010110101010",
				"011010101011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110011010",
				"010010011010",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011010111011",
				"011110111100",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"011110111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010101110111",
				"001101010101",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110011",
				"001000110011",
				"001101000100",
				"001101100101",
				"010001110110",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110111011",
				"100010111100",
				"100111001100",
				"100010111100",
				"100010111011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001110111",
				"010001110111",
				"010101110111",
				"011010001000",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010101111000",
				"010010001000",
				"010010001000",
				"001110001000",
				"001110000111",
				"010001110111",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100111",
				"010101100111",
				"010101100111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101010110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101100101",
				"001101100110",
				"001101100111",
				"011110111100",
				"100111011110",
				"100111101111",
				"100111101111",
				"011111011101",
				"100011101110",
				"100011011110",
				"011111011110",
				"100011011111",
				"100011011110",
				"011111011110",
				"100011101111",
				"100011011111",
				"011111011111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100111011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101111111111",
				"101111101111",
				"101011011101",
				"011110011001",
				"010101010101",
				"001100110011",
				"010001000100",
				"010101010110",
				"100110011011",
				"101111001101",
				"110111101111",
				"101111001101",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010101010",
				"100110000111",
				"100001010100",
				"100101010100",
				"100101010100",
				"100101010100",
				"100101010100",
				"011101010100",
				"011101100110",
				"011110001001",
				"100110101100",
				"100011001110",
				"011111001110",
				"011011001110",
				"011011001110",
				"100011001111",
				"100111011111",
				"101011011111",
				"101011101111",
				"101011111111",
				"101011101111",
				"100111011110",
				"100011001110",
				"100011001110",
				"011111001101",
				"011011001101",
				"011011001101",
				"010111001101",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111101",
				"011010111100",
				"010110101100",
				"010110101100",
				"010110111100",
				"011010111100",
				"010110101100",
				"010010101011",
				"010110101011",
				"011010111101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011110111101",
				"100011001101",
				"100010111101",
				"011110101011",
				"011110011011",
				"011110011011",
				"011010011011",
				"010110011100",
				"010010011100",
				"010110101101",
				"011010101101",
				"011010011100",
				"100010101100",
				"100010011100",
				"011101111001",
				"100001100110",
				"100001100101",
				"100101100101",
				"100101010100",
				"100001000010",
				"011000100001",
				"011000110010",
				"011101100101",
				"100110011001",
				"100110111100",
				"100111001101",
				"100011001101",
				"011110111101",
				"011111001110",
				"100011001110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"100011001100",
				"100011011100",
				"100111011101",
				"100111011101",
				"101011011101",
				"101111011110",
				"101111011101",
				"101011001101",
				"101011001101",
				"101011011100",
				"101011011100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111001100",
				"101111001101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101111001100",
				"101111011100",
				"101011011100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011011101",
				"100111011101",
				"100111001101",
				"011111001100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111011",
				"011010111011",
				"010110101010",
				"010110011010",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"010110011011",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010001100110",
				"001101010101",
				"000100110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100010",
				"001100110100",
				"010001010101",
				"010101100110",
				"011001110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110101010",
				"011110101010",
				"011110111010",
				"011110111011",
				"011110111011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110101011",
				"100010101011",
				"011110011011",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110101011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100110",
				"011110101011",
				"101111111111",
				"100111101110",
				"101011101111",
				"100011011101",
				"100111101110",
				"100111101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111101111",
				"101111101110",
				"110011101110",
				"101111001100",
				"100110101010",
				"100010011001",
				"100110111011",
				"101111011101",
				"101111101110",
				"110011101111",
				"110011111111",
				"101111011110",
				"101111001101",
				"101010111011",
				"101110111011",
				"110010101010",
				"101010000111",
				"100001010100",
				"100101010100",
				"100101010100",
				"100101010100",
				"100101010100",
				"100001100101",
				"100001100111",
				"011101111000",
				"100110101011",
				"100111001110",
				"100011001111",
				"011010111110",
				"010110111101",
				"011110111101",
				"100111001111",
				"101011011111",
				"101011011111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111001110",
				"011111001101",
				"011111011110",
				"011011001101",
				"011011001101",
				"011010111101",
				"100011001110",
				"100111011111",
				"011111001101",
				"011111011110",
				"011111001101",
				"011011001101",
				"011010111100",
				"010110101100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101100",
				"010110101100",
				"010110101100",
				"011010111101",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011110111101",
				"011110101100",
				"011110011010",
				"011110011011",
				"011110011011",
				"011010011011",
				"010110001011",
				"010010001011",
				"010110101101",
				"011010101101",
				"011010011100",
				"011110101100",
				"100110101100",
				"100110011010",
				"100101111000",
				"100001010101",
				"100001010100",
				"100101010101",
				"100001000011",
				"011000100010",
				"011000110011",
				"100001100110",
				"101010101011",
				"101010111100",
				"100110111101",
				"100010111110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101111011101",
				"101011001101",
				"101111001101",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011101110",
				"110011101110",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001100",
				"101011001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011011100",
				"101011001100",
				"101011011101",
				"101011011101",
				"101011011101",
				"100111001100",
				"011111001100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110011010",
				"010110101011",
				"011010101011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010010011010",
				"010110011010",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110101011",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110001001",
				"010001111000",
				"010001100110",
				"001101010101",
				"001000110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110011",
				"010001010101",
				"010101110111",
				"011010001000",
				"011110011001",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110011010",
				"011110011011",
				"011110101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010101100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"011010011010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"010001100110",
				"010001110111",
				"010001100110",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100110",
				"011010011010",
				"101111111111",
				"101111101111",
				"101111111111",
				"100111011110",
				"101011101110",
				"101011111111",
				"100111101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011101110",
				"110011101110",
				"110011101110",
				"110011101110",
				"110011111110",
				"110011111111",
				"101111101110",
				"101111111111",
				"101111101111",
				"110011101111",
				"110011011110",
				"101110111100",
				"110010101011",
				"101110011001",
				"100101110110",
				"100001010100",
				"100101010100",
				"101001010100",
				"101001010100",
				"101001100101",
				"100101110110",
				"101010001000",
				"100110001001",
				"100110101011",
				"101011001110",
				"100111011111",
				"100011011111",
				"011010111101",
				"011010101101",
				"100011001110",
				"100111011111",
				"100111001111",
				"100011011111",
				"100011011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100011011110",
				"011111001110",
				"011011001101",
				"011010111101",
				"011110111101",
				"100111011111",
				"100111011111",
				"011010111101",
				"011011001101",
				"011010111101",
				"010110111100",
				"010110111100",
				"010110101011",
				"010110101011",
				"010010011011",
				"010010011010",
				"010010011010",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110011011",
				"011110011010",
				"100010011011",
				"100010011011",
				"011110011011",
				"010110001010",
				"010110001011",
				"010110011100",
				"011010011100",
				"011010011011",
				"011110011011",
				"100010101100",
				"101010101100",
				"101010011010",
				"100101111000",
				"011101010101",
				"011101000100",
				"011101000100",
				"011000110011",
				"011001000100",
				"100110001001",
				"101110111101",
				"101010111101",
				"100010111101",
				"100010111110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101111011100",
				"101011001100",
				"101011001100",
				"101011011101",
				"100111011101",
				"100011001100",
				"011110111100",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010010011001",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101010",
				"010010011010",
				"010010101010",
				"010110101011",
				"010110111011",
				"011010111011",
				"010110111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111011",
				"011010111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110101011",
				"010110011001",
				"010110011001",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001000",
				"010101111000",
				"010001110111",
				"001101010101",
				"001000110011",
				"000000100010",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000100010",
				"001001000100",
				"001101010101",
				"010101110111",
				"011010001000",
				"010110001000",
				"011010011001",
				"011110101010",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011110101011",
				"011110101011",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010101100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111100",
				"100010111100",
				"100110111101",
				"101010111101",
				"101010111101",
				"100110101100",
				"100110101100",
				"100010111100",
				"100010111100",
				"011110111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010001001",
				"010101111000",
				"010110001001",
				"011010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100110",
				"011010001001",
				"101111101110",
				"110111111111",
				"110011111111",
				"101111101111",
				"101011011101",
				"101111111111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100011101110",
				"100011101111",
				"100111101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101110",
				"110011101110",
				"110011111110",
				"110011111110",
				"101111111110",
				"101011111110",
				"101011111110",
				"101111111111",
				"101111101111",
				"110111111111",
				"110111101111",
				"110111011110",
				"110110111100",
				"101110011001",
				"100001100110",
				"100001010100",
				"101001010100",
				"101001100101",
				"101001100100",
				"101001100101",
				"100101100101",
				"100101110111",
				"101010001001",
				"101010101011",
				"101011001101",
				"101011011111",
				"100111011111",
				"011111001110",
				"011110111101",
				"100010111110",
				"101011011111",
				"100111001111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111011111",
				"011111001110",
				"011010111101",
				"010110101011",
				"011110111101",
				"100111011111",
				"011110111101",
				"011010111101",
				"011011001101",
				"010110111100",
				"010110111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010010101011",
				"010010011010",
				"010010011010",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011010111100",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010101011",
				"011010011010",
				"100010011010",
				"100110101011",
				"100010011011",
				"011110001010",
				"011010001010",
				"010110001011",
				"010110011011",
				"010110011011",
				"010110011011",
				"011010011011",
				"100010101100",
				"100110101100",
				"101010111100",
				"101110101100",
				"100110001001",
				"011101010110",
				"011001000100",
				"010100110100",
				"100001100111",
				"101110111100",
				"101111001101",
				"100110111101",
				"100010111101",
				"100011001110",
				"100011001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100111001101",
				"100111001101",
				"101011001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111011100",
				"101111011100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111011100",
				"100011001100",
				"011111001100",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110011011",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110101011",
				"010110011010",
				"010110101010",
				"011010111011",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001110111",
				"001101010110",
				"001001000100",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"000100110011",
				"001001000101",
				"010001100110",
				"010101111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011110111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110101011",
				"100010101100",
				"100110111100",
				"101010111101",
				"101010111101",
				"100110101100",
				"100110101100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110001001",
				"010101111000",
				"010101111000",
				"011010001001",
				"011110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010001001",
				"010101111000",
				"010101110111",
				"010101111000",
				"010110001000",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101100110",
				"001101100101",
				"001101100101",
				"001101100110",
				"001101010101",
				"010101110111",
				"101011001100",
				"111011111111",
				"110111111111",
				"110011111111",
				"101011011101",
				"101111101110",
				"101011111111",
				"101011111111",
				"101011101111",
				"100011011110",
				"011111001101",
				"100011011110",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111110",
				"110011111110",
				"101111111111",
				"101111111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110111101111",
				"111011101111",
				"111011011110",
				"111011001100",
				"101010001000",
				"100101100101",
				"100101010100",
				"100101010100",
				"101001010100",
				"101001100101",
				"100101100101",
				"100101110110",
				"100001110111",
				"101010101011",
				"101111001110",
				"101011011111",
				"100111011111",
				"100111011111",
				"100010111110",
				"100010111101",
				"100111001111",
				"100111001110",
				"100011001110",
				"100011011110",
				"011111011110",
				"100011011111",
				"100011101111",
				"100011011111",
				"011111001110",
				"011010111100",
				"011010101011",
				"100111011110",
				"100111011111",
				"011110111101",
				"011011001101",
				"011011001101",
				"010110111100",
				"010110111100",
				"010110101011",
				"010110101011",
				"010010101011",
				"010010101011",
				"010110101011",
				"010110101011",
				"010110011011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011010111100",
				"011010101010",
				"011010011010",
				"100010101010",
				"100110101011",
				"100010011010",
				"011110001001",
				"011110001010",
				"011010011011",
				"010110011011",
				"010110011011",
				"011010011011",
				"011110101100",
				"011110101100",
				"100010101100",
				"100110111101",
				"101010111101",
				"101110111101",
				"101010011011",
				"011101100111",
				"100001111000",
				"101010101011",
				"101111001101",
				"101011001101",
				"100111001101",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100111001101",
				"100111001101",
				"101011001101",
				"101111001101",
				"110011001110",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"100111001101",
				"101011001101",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100111001100",
				"100011001100",
				"011110111011",
				"011010111011",
				"010110101010",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011010101010",
				"011010111011",
				"011111001100",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010111001100",
				"010111001100",
				"010111001100",
				"010111001100",
				"010111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101100",
				"011010111011",
				"011010111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010101111000",
				"010001100110",
				"001001000011",
				"000000100001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000100010",
				"000100110011",
				"001101010101",
				"010001110111",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011110111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111101",
				"100010111100",
				"011110101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010111011",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"100010101100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110101100",
				"100110101100",
				"100010101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110101010",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011010001001",
				"010101111000",
				"010101111000",
				"011010001001",
				"011110101010",
				"011110101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010001001",
				"010101111000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101110110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001110110",
				"010001110110",
				"001101100110",
				"010101110111",
				"100010111011",
				"110111111111",
				"110111111111",
				"110111111111",
				"101111101110",
				"101111101110",
				"110011111111",
				"110011111111",
				"101111101111",
				"101011011110",
				"100011001100",
				"100011001101",
				"101011011110",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101110",
				"110011101111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110011101110",
				"110011111110",
				"110011111110",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011101111",
				"110011101110",
				"111011111111",
				"111011101111",
				"111111111111",
				"111011011100",
				"101010011000",
				"100101100101",
				"100001000100",
				"100101010100",
				"101001110110",
				"101001110110",
				"100101110111",
				"101010001000",
				"110010111100",
				"110011011111",
				"101111011111",
				"101011011111",
				"101011011111",
				"100111001110",
				"011110101101",
				"100010111110",
				"100010111110",
				"011110111110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"010110101011",
				"011110111101",
				"101011101111",
				"100111011111",
				"011010111101",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010010101100",
				"010010101011",
				"010010101011",
				"010010011011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"011010011010",
				"011110011010",
				"100110101011",
				"100110101011",
				"100010011010",
				"011110001010",
				"011110001010",
				"011010011010",
				"011010011011",
				"010110011011",
				"011010011100",
				"011110101100",
				"011110101100",
				"100010101101",
				"100010101101",
				"100010101100",
				"100110111101",
				"101111001110",
				"101010111100",
				"101010111100",
				"101111001101",
				"101011001101",
				"100111001101",
				"100011001101",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011001101",
				"100111001101",
				"101011001101",
				"101111011101",
				"110011011110",
				"110011001110",
				"110011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100011001101",
				"100111001101",
				"101011011101",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111011100",
				"100111001100",
				"100011001100",
				"011010111011",
				"011010101010",
				"010110101010",
				"011010101011",
				"010110101010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"010111001100",
				"010111001100",
				"010110111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010011011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010101110111",
				"010001100110",
				"001001000011",
				"000000100001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"001001000100",
				"010001100110",
				"010001110111",
				"010110001000",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111011",
				"011010101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011010011011",
				"011010011011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"011110101011",
				"011010011010",
				"011010011010",
				"011110101011",
				"100010111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100110111101",
				"100111001101",
				"100110111101",
				"100010101100",
				"100010101100",
				"100010101100",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010011010",
				"011110011010",
				"011110011010",
				"011010001001",
				"010101111000",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"011010001001",
				"011110001001",
				"011110001001",
				"010101110111",
				"010001100110",
				"010101110111",
				"011010001001",
				"011010001001",
				"010101111000",
				"010001110111",
				"010001110111",
				"010010001000",
				"010010001000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110110",
				"001101110110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101111000",
				"100010101011",
				"110011101111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101111",
				"101011011110",
				"101011011101",
				"101111011110",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101110",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"101111011110",
				"110111111111",
				"110111101110",
				"111111111111",
				"111111111111",
				"110010111010",
				"101001110111",
				"100101010101",
				"100101100101",
				"101001110110",
				"100101110110",
				"100101110111",
				"110010111011",
				"110111011110",
				"110111101111",
				"101111011111",
				"101011011111",
				"100111011111",
				"100010111110",
				"011110011101",
				"100110111110",
				"100010101101",
				"011110111101",
				"011110111101",
				"011011001101",
				"011011001110",
				"011011001110",
				"011010111101",
				"011111001110",
				"010110101100",
				"100011001110",
				"101011101111",
				"100011011110",
				"011011001101",
				"010110111100",
				"010111001100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010010101011",
				"010010101011",
				"010010101011",
				"010110101011",
				"011010101100",
				"011010111100",
				"011110111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110101011",
				"100110101100",
				"100110101011",
				"100010011010",
				"100010011010",
				"011110001010",
				"011110011011",
				"010110001010",
				"010110001011",
				"011010011100",
				"011110101101",
				"100010111101",
				"100010111110",
				"011110111101",
				"011110101100",
				"011110101100",
				"100111001110",
				"101111011111",
				"101011011110",
				"100111001101",
				"100111001101",
				"100111001110",
				"100011001101",
				"011111001110",
				"011111001101",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100111011101",
				"101111011101",
				"101111011110",
				"110011011110",
				"110011011110",
				"101111001101",
				"101011001100",
				"100111001101",
				"100111011101",
				"100111011101",
				"100011011101",
				"100111011101",
				"101011011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"101111001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111011100",
				"101111011101",
				"101111011100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011011101",
				"100111001100",
				"011110111011",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"010110011010",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110101010",
				"011010111011",
				"011010111011",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101010",
				"010010011010",
				"010010011001",
				"010010011001",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011011",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011001",
				"010110001000",
				"010101110111",
				"001101010101",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100010",
				"001001000100",
				"010001100110",
				"010101111000",
				"011010011001",
				"011010011001",
				"011110101010",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"100011001101",
				"011110111100",
				"011010101011",
				"011110101011",
				"100010111100",
				"100110111101",
				"100010101100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011011001100",
				"010111001100",
				"010111001100",
				"010111001100",
				"010110111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110111100",
				"011110111011",
				"011110111100",
				"011110111100",
				"100011001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011011001100",
				"011010111011",
				"011110111100",
				"100010111100",
				"011110101011",
				"011110101011",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"010110101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"011001111001",
				"011001111000",
				"010001100111",
				"001101010110",
				"010001010110",
				"010101111000",
				"011010001000",
				"010101111000",
				"010101111000",
				"010110001001",
				"001101110111",
				"010001110111",
				"010010001000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110110",
				"001101110110",
				"001101110111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001110111",
				"010101111000",
				"010101111000",
				"100110111100",
				"101111101111",
				"101111011110",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"101111101110",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101110",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011101110",
				"110011111111",
				"110111111111",
				"111111111111",
				"111111101110",
				"110110111011",
				"101010001000",
				"100001100101",
				"100001100110",
				"101010011000",
				"110011001100",
				"111111101111",
				"111011101111",
				"110111101111",
				"101111011111",
				"101011011111",
				"101011011111",
				"100111001111",
				"100010111110",
				"100110111110",
				"100110111110",
				"100011001110",
				"011111001110",
				"011111001110",
				"011011001110",
				"011011001110",
				"011111001110",
				"011010111101",
				"011010111100",
				"100011011110",
				"100011011111",
				"011111001101",
				"011011001101",
				"010110111100",
				"010111001101",
				"010111001100",
				"010110111101",
				"010110111100",
				"010110111100",
				"010110101100",
				"010110101011",
				"010110101011",
				"010110101100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010101100",
				"010110101011",
				"011010101100",
				"010010011011",
				"010110101011",
				"011110101100",
				"100010101100",
				"100010101011",
				"100110101011",
				"100110011011",
				"100010011011",
				"011110011011",
				"011110011011",
				"011010011011",
				"011010011100",
				"011010011100",
				"011110111110",
				"011110111110",
				"011110111110",
				"011110111110",
				"011110111101",
				"100010111101",
				"100111001110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011101",
				"100111011101",
				"101011011101",
				"110011011110",
				"110011011110",
				"110011011101",
				"101111001101",
				"101011001100",
				"100111001100",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100111011101",
				"101011011101",
				"101111001101",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011001100",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011011100",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100111011100",
				"100011001100",
				"011110111011",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"001110001000",
				"010010011001",
				"011010101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"010110101011",
				"010010011010",
				"010010011001",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111011",
				"011111001100",
				"011111001100",
				"011010111100",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011011001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010110001001",
				"010110001000",
				"010001100110",
				"000101000011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100110011",
				"001101010101",
				"010101110111",
				"011010001001",
				"011110011010",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011010101100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011111001100",
				"011110111100",
				"011110101011",
				"011110101011",
				"100010111100",
				"100110111101",
				"100010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"010111001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011110111100",
				"011110111100",
				"011110101100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011011001100",
				"011010111011",
				"011110111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"011110111011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"001110001000",
				"001101111000",
				"010001111000",
				"010110001001",
				"011010001001",
				"011110001001",
				"011001111000",
				"010101110111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"010001100111",
				"010001100111",
				"010001111000",
				"010001111000",
				"011110101011",
				"101011011110",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111110",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101110",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111101110",
				"111111111111",
				"111111111111",
				"111011001100",
				"101110101010",
				"101110101010",
				"110111001100",
				"111111111111",
				"111111111111",
				"111011101111",
				"110011101111",
				"101011011111",
				"100111011111",
				"100111011111",
				"100111001111",
				"100110111110",
				"101011001111",
				"101011001111",
				"100111001110",
				"011110111110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011010111101",
				"100011001110",
				"100111101111",
				"100011011110",
				"011011001101",
				"011011011101",
				"011011011101",
				"010111001101",
				"010111001101",
				"010110111101",
				"010110111100",
				"010110111100",
				"010110101100",
				"010110101100",
				"010110101100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111101",
				"011110111101",
				"011110111101",
				"011010111100",
				"010110101011",
				"010110101011",
				"011010101100",
				"011110111100",
				"100010111100",
				"100010101100",
				"100010011011",
				"100010011011",
				"011110001010",
				"011110011011",
				"011110011100",
				"011010011011",
				"011010011100",
				"011010101100",
				"011110111110",
				"011110111110",
				"011110111110",
				"011110111101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111011101",
				"100111011101",
				"101011011101",
				"101111011110",
				"110011011110",
				"110011011101",
				"101111001101",
				"101011001100",
				"100111001100",
				"100011001101",
				"100011011101",
				"100111011110",
				"100111011101",
				"100111011101",
				"101011011101",
				"101111011101",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011011100",
				"110011011101",
				"110011011101",
				"110011011100",
				"101111001100",
				"101111011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"101011001101",
				"100111011101",
				"100111001100",
				"100011001100",
				"011110111011",
				"011010101010",
				"010110011001",
				"010010011001",
				"010010001001",
				"001110001000",
				"001110001000",
				"010010011001",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010010011010",
				"010010011001",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111011101",
				"011111001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010001110111",
				"001001010101",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000000100010",
				"001001000100",
				"001101010110",
				"010110001000",
				"011110011001",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110111011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011010111101",
				"011010111101",
				"011110111101",
				"100010111101",
				"100111001110",
				"100011001101",
				"011110111100",
				"011010101100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011111001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100110111101",
				"100010111101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011110111100",
				"011110111100",
				"100010101100",
				"100110111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010011010",
				"011110011010",
				"011010011011",
				"011010101011",
				"011010111011",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010110001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001001",
				"010110001000",
				"010101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101100111",
				"010001111000",
				"010001111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001101000",
				"010001100111",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001111000",
				"010001111000",
				"011010011010",
				"101011001110",
				"110011101111",
				"101111011110",
				"101111101110",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101110",
				"111011101111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111111101111",
				"111111101111",
				"111111101111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101111",
				"101011011111",
				"100111011111",
				"100111011111",
				"100111001111",
				"100111001111",
				"101011001111",
				"101011001111",
				"100111001110",
				"100010111110",
				"100011001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"100111101111",
				"100111101111",
				"011111001110",
				"011011001101",
				"011011011101",
				"011011011101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"100011001110",
				"011111001101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011010111100",
				"010110011011",
				"010110011011",
				"011010101100",
				"011110101100",
				"011110101100",
				"011110011011",
				"011110011011",
				"011110011011",
				"011010001010",
				"011010011011",
				"011010011011",
				"010110011011",
				"010110011100",
				"011010101100",
				"011110111110",
				"011110111110",
				"011110111101",
				"011110111101",
				"100011001110",
				"100111001110",
				"100011001110",
				"100111001110",
				"101011001110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011101",
				"100111001101",
				"100111011110",
				"101011011110",
				"100111011101",
				"101011011101",
				"101011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111001101",
				"101011001100",
				"100111001100",
				"100011001100",
				"100111011101",
				"100111011110",
				"101011011101",
				"101011011101",
				"101111011101",
				"101111011101",
				"101111001100",
				"110011011101",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011101",
				"110011011101",
				"110011011100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001100",
				"100111001100",
				"100111001100",
				"100011001100",
				"011110111100",
				"011110111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010010011001",
				"010010011010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010011011",
				"011010011011",
				"011110101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001000",
				"001101100110",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001001000100",
				"010001010110",
				"010001110111",
				"011010001000",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011110111101",
				"100010111101",
				"100111001110",
				"100111001110",
				"100010111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"100010111100",
				"100011001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100110111101",
				"100010111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010101010",
				"011010011010",
				"011110001010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"011010011001",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010101111000",
				"010101111000",
				"010101111000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010101111000",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"001101100111",
				"001001010110",
				"001101100111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010001101000",
				"010001111000",
				"010001100111",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001111000",
				"010110001001",
				"010110001001",
				"100111001101",
				"110111111111",
				"110011101111",
				"101111011110",
				"101111011101",
				"101111101110",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101110",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110011011111",
				"101111011111",
				"101011011110",
				"100111011110",
				"100111011111",
				"100111001111",
				"101011001111",
				"101011001111",
				"101011001110",
				"100110111110",
				"100110111110",
				"100111011110",
				"100011011110",
				"011111001110",
				"011111001101",
				"100111011111",
				"101011101111",
				"100011011110",
				"100011011110",
				"100011101110",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011010101100",
				"010110011010",
				"011010011011",
				"011010011100",
				"010110001010",
				"011010001010",
				"011110011100",
				"011110101100",
				"011010001011",
				"011010011011",
				"010110011011",
				"010110011011",
				"010110011100",
				"011010101101",
				"011110111110",
				"011110111110",
				"011010101101",
				"011110111101",
				"100010111101",
				"100011001110",
				"100010111110",
				"100111001110",
				"100111001110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011011101",
				"101111011101",
				"101111011101",
				"110011011110",
				"110011011110",
				"110011011101",
				"101111001101",
				"101011001101",
				"100111001100",
				"100111001101",
				"101011011110",
				"101011011101",
				"101011001101",
				"101111011101",
				"110011011101",
				"110011001100",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011011100",
				"110111011101",
				"110011011101",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110101100",
				"011110101011",
				"011010011011",
				"011010011011",
				"011110101011",
				"011110101100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010011010",
				"010110001001",
				"011010011010",
				"011010011011",
				"011110101011",
				"011110101100",
				"011010101100",
				"011010101100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010001111000",
				"001101100110",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000100010",
				"001101010101",
				"010101110111",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100010111101",
				"100110111110",
				"100111001110",
				"100110111101",
				"100011001101",
				"100111001110",
				"100011001110",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011011001100",
				"011111001101",
				"100011001101",
				"100111001101",
				"100110111100",
				"100010101100",
				"100010101011",
				"100110111100",
				"100111001101",
				"100111001100",
				"100010111100",
				"011110101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010011010",
				"011110001001",
				"011001111000",
				"010101100111",
				"010101100111",
				"010101100111",
				"010101111000",
				"010110001001",
				"011010101010",
				"011110101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"011010011010",
				"010110011001",
				"011010011001",
				"011010001001",
				"010101111000",
				"010001100111",
				"010001010111",
				"010001100111",
				"010001110111",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"001101100111",
				"001101100110",
				"001101010110",
				"001101100110",
				"010001110111",
				"011010001000",
				"011010001000",
				"011001111000",
				"010101111000",
				"010001110111",
				"001101100111",
				"001101100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010101111000",
				"001101100111",
				"011010011010",
				"101111101111",
				"110111111111",
				"110111111111",
				"101111101110",
				"101111011101",
				"110011101110",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011101111",
				"110111101111",
				"110111111111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101111011111",
				"100111011110",
				"100111011110",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011001110",
				"100110111101",
				"100010111101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"101111111111",
				"101111101111",
				"100011011110",
				"100111011111",
				"100111101111",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011010101100",
				"011010101100",
				"011010011100",
				"011010011011",
				"011010011100",
				"011110101101",
				"011110101101",
				"011010011100",
				"010110011100",
				"010110011011",
				"010110101100",
				"010110101100",
				"011010111101",
				"011110111110",
				"011110111110",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"100010111110",
				"100011001110",
				"100111001110",
				"100111001110",
				"101011011110",
				"101011011111",
				"100111011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001110",
				"101011001101",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"101111011101",
				"101011001101",
				"101011001100",
				"101011001101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011011101",
				"110011011101",
				"101111001100",
				"101111001100",
				"101111011101",
				"101011011101",
				"101011011101",
				"100111001100",
				"100011001100",
				"100011001100",
				"100111001101",
				"100011001100",
				"011110111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"010111001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010011011",
				"011110101011",
				"011110101100",
				"011110111101",
				"011110111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010011010",
				"010110001001",
				"011010011010",
				"011110101011",
				"011110101100",
				"011110101100",
				"011010101100",
				"011010101100",
				"010110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010010001001",
				"010001110111",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101010101",
				"010110001000",
				"011010011001",
				"011110101010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011110111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100111001110",
				"100110111110",
				"100110111101",
				"100010111101",
				"100011001110",
				"100111011110",
				"100011001110",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011110",
				"100011011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011111001101",
				"100010111101",
				"100110111100",
				"100110011011",
				"100010001010",
				"100010001010",
				"100110101011",
				"100110111100",
				"100010111011",
				"011010101010",
				"011010101011",
				"011010111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011011001100",
				"011110111011",
				"011110111011",
				"100010011010",
				"011001111000",
				"010101010110",
				"010101010110",
				"011001100111",
				"011110001001",
				"011110101010",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110001001",
				"010101100111",
				"010101010110",
				"010101100111",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010001111000",
				"010001110111",
				"001101100111",
				"001101010110",
				"010001100110",
				"010001100111",
				"010101100111",
				"010001100111",
				"010001100111",
				"001101100111",
				"001101100110",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001111000",
				"001101100111",
				"010001100111",
				"011110101010",
				"101111101110",
				"111011111111",
				"110111111111",
				"110111111110",
				"110111101110",
				"110111101110",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101110",
				"110111101110",
				"111011111111",
				"111111111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011111111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011111",
				"101011011110",
				"100111101111",
				"101011101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"101011011111",
				"100110111101",
				"100010111100",
				"100010111101",
				"100011001101",
				"100111011110",
				"101011101111",
				"101111101111",
				"101011101111",
				"100111011110",
				"100111011110",
				"100111011111",
				"100011011110",
				"100111001110",
				"100010111101",
				"100011001100",
				"100111001101",
				"100111001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100111001101",
				"100010111100",
				"100111001101",
				"100010111101",
				"100010111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111101",
				"011110101100",
				"011110101100",
				"100010111101",
				"100010111110",
				"011110101101",
				"011010101101",
				"011010101101",
				"010110101100",
				"010110101100",
				"010110111100",
				"010110111101",
				"011010111101",
				"011110111101",
				"011110111110",
				"011110111101",
				"011111001110",
				"011110111101",
				"011110111101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111011110",
				"101011011111",
				"100111011110",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001110",
				"100111001110",
				"100111001101",
				"101011011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001101",
				"101011001100",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110111011101",
				"110111011101",
				"110011011100",
				"110011011100",
				"110011011101",
				"101111001100",
				"101111001100",
				"101111011101",
				"101011011101",
				"101011011101",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011010111011",
				"010110101010",
				"010010011010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101010",
				"010110101010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011010111011",
				"011010111011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011010111011",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"011111011101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100011001100",
				"100011001100",
				"100011001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111011",
				"011110101100",
				"011110111100",
				"100010111101",
				"100010111101",
				"100011001101",
				"011110111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"100010111100",
				"011110101011",
				"011110011010",
				"011010001001",
				"011010011010",
				"011110101011",
				"011110101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101010",
				"010110101010",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001000",
				"001101010101",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100110011",
				"001101010101",
				"010101111000",
				"011010011001",
				"011110011010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011111001101",
				"100011001101",
				"100111001101",
				"101110111101",
				"101110101100",
				"101010011011",
				"101110101011",
				"101010111100",
				"100110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100010101011",
				"011101111000",
				"011001010110",
				"011101010111",
				"100110001001",
				"100110101011",
				"100010111100",
				"011010111011",
				"010110111010",
				"010110101010",
				"011010101011",
				"011110111011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110001001",
				"011001100111",
				"011001100111",
				"011101111000",
				"011110001001",
				"011110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011000",
				"010010011000",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010110001001",
				"010110001000",
				"010101111000",
				"010001100111",
				"010001010110",
				"001101010101",
				"001101000101",
				"001101010110",
				"001101100110",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"001101100111",
				"010001100111",
				"001101010110",
				"010001100111",
				"101011001100",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101110",
				"110111101110",
				"111011111111",
				"111111111111",
				"111011111111",
				"110111011110",
				"110111101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111110",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101110",
				"111011111111",
				"111011111111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011001110",
				"101011001110",
				"101011011110",
				"101011101111",
				"101111111111",
				"101111011111",
				"101011011110",
				"100111011110",
				"100011001110",
				"100011001101",
				"100111001110",
				"100110111101",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001110",
				"100111011110",
				"100111001101",
				"100011001101",
				"100010111101",
				"011110101100",
				"011110101100",
				"100011001110",
				"100011001110",
				"011110111110",
				"011110111110",
				"011010111110",
				"010110111101",
				"010110111101",
				"011011001101",
				"011010111101",
				"011111001110",
				"011110111101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011011110",
				"100111011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"101011001101",
				"101011011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101011001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110111011101",
				"110111011101",
				"110011011100",
				"110011011101",
				"110011011101",
				"101111001100",
				"101011001100",
				"101011011101",
				"101011011101",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011111001100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010010101010",
				"010010101010",
				"010010101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"011111011110",
				"011111011101",
				"011011011101",
				"011011001100",
				"011011001100",
				"011011001011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100011001011",
				"100011001100",
				"100011001100",
				"100011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001101",
				"011111001100",
				"011111001100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"011010011010",
				"011010011010",
				"011110101011",
				"011110111100",
				"011110111100",
				"011010111101",
				"011010111101",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011011",
				"010110011010",
				"010110001001",
				"010001100110",
				"001000110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100110011",
				"010001100110",
				"010110001000",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010111011",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001110",
				"100111001101",
				"100010111101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011011110",
				"011111001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100110111100",
				"100110111100",
				"100010101011",
				"100110111100",
				"100110111100",
				"100010111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011011001101",
				"011011001101",
				"010111001101",
				"011011001101",
				"011111011101",
				"100011001101",
				"101011001101",
				"110010111101",
				"101110101100",
				"110010101100",
				"110010111101",
				"101110111100",
				"100010101011",
				"011010111010",
				"011011001011",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110101010",
				"010101110111",
				"010101000110",
				"011101100111",
				"100110001010",
				"100110101011",
				"100010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"011010101010",
				"011110101010",
				"011110001001",
				"010101100111",
				"011001100111",
				"011110001001",
				"100010011010",
				"011110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011000",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101100111",
				"010001010110",
				"001001000100",
				"001001010101",
				"001101100111",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"001101100111",
				"001001010110",
				"010001100111",
				"001101010110",
				"010001110111",
				"101111011101",
				"111011111111",
				"110111111111",
				"111011111111",
				"111111111111",
				"111011101111",
				"111011101110",
				"111011101111",
				"111111111111",
				"111011111111",
				"110111101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110011011110",
				"101111011110",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"110011111111",
				"101111101111",
				"100111001101",
				"101011011110",
				"100111001101",
				"100011001101",
				"100111001101",
				"100110111101",
				"101010111101",
				"101010111100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101010111100",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011001101",
				"100111001101",
				"101011011110",
				"100111001101",
				"100111001101",
				"100110111101",
				"100110111101",
				"100110111101",
				"100110111110",
				"100010111110",
				"100011001110",
				"100011001110",
				"011111001110",
				"011010111101",
				"010111001101",
				"011011011110",
				"011011001101",
				"011111011110",
				"011011001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011101110",
				"100011011110",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"101011001101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011101",
				"110111011101",
				"110011011101",
				"110011011100",
				"110011011101",
				"110011011100",
				"101111001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010101010",
				"010010011001",
				"010010011001",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"010010101010",
				"010010011010",
				"010010101010",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110101011",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011011001100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111011",
				"011110111011",
				"100010111100",
				"100011001100",
				"100011001100",
				"011111001100",
				"011110111011",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"011111001110",
				"011111001110",
				"011011001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"011110101100",
				"011010011010",
				"011010011011",
				"011010101011",
				"011010101100",
				"011110111101",
				"011011001101",
				"011010111101",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101011",
				"010110011011",
				"010110011010",
				"010101110111",
				"001101000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000100110011",
				"010001100110",
				"010110011000",
				"011010101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100111001110",
				"100110111101",
				"100110111101",
				"100010111101",
				"100010111100",
				"100010111101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"100011001101",
				"100110111100",
				"100110101011",
				"100010011010",
				"011101111001",
				"100110011010",
				"101010101011",
				"100110111100",
				"100010111011",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011011001101",
				"011011001101",
				"011111011110",
				"011011001101",
				"011011001101",
				"011111011101",
				"011111011110",
				"100011001101",
				"100111001101",
				"101011001101",
				"101110111101",
				"101110111101",
				"101110101100",
				"101010101100",
				"100110101100",
				"100010111011",
				"011111001100",
				"011111011100",
				"011111011101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010101010",
				"011010001001",
				"011001111000",
				"010101111000",
				"011110011010",
				"100010101011",
				"100010111100",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110111010",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111010",
				"010110101010",
				"010110111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110001000",
				"010001100111",
				"010001100111",
				"010101101000",
				"011010001001",
				"011110101011",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010101111000",
				"010101111000",
				"010001100111",
				"010001010110",
				"001101000101",
				"010101110111",
				"011010001000",
				"010110001000",
				"010001110111",
				"010101110111",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"001101100110",
				"010001110111",
				"010110000111",
				"101111011101",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101110",
				"111011111111",
				"110111101110",
				"111011101110",
				"111011101110",
				"110111101110",
				"110111101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"111011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110011101110",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101110",
				"110011101111",
				"110011111111",
				"101111101110",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"110011101111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110011101110",
				"101111011110",
				"101111011110",
				"101011011101",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001101",
				"101011001101",
				"101111001101",
				"101010111100",
				"110011011101",
				"110111101110",
				"110011001101",
				"101111001101",
				"110011011110",
				"101111001101",
				"110011011110",
				"101111001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101010111101",
				"101111001101",
				"101010111101",
				"100111001101",
				"101011001110",
				"100011001110",
				"100011001110",
				"011111011110",
				"011011001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001100",
				"110011001100",
				"110011011101",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011011100",
				"110011011101",
				"101111011100",
				"101111001100",
				"101011001100",
				"100111001100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001100",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110111010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011010111011",
				"010110101010",
				"010110101011",
				"011010111100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100010111100",
				"100010111100",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011011001100",
				"010111001100",
				"010111001100",
				"010111001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001110",
				"011011001110",
				"011011001101",
				"011011001110",
				"011011001110",
				"011011001101",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111101",
				"011110111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011001",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110001000",
				"001101010110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"010001100110",
				"010110001000",
				"011010101010",
				"011010111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"100111001110",
				"100110111110",
				"100110111101",
				"100111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"010111011101",
				"011011011101",
				"011011011101",
				"100011011110",
				"100111001101",
				"101010111100",
				"100110101011",
				"100110001010",
				"100010001001",
				"101010101011",
				"101111001100",
				"101011001101",
				"100111001100",
				"011111001100",
				"011111011101",
				"011011011100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"101010111101",
				"101111001101",
				"101010111101",
				"101010111101",
				"100110111100",
				"100110111100",
				"100011001100",
				"011111001100",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101010",
				"011010101010",
				"011110111011",
				"100010111100",
				"100010111100",
				"011110111011",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"010110001001",
				"011010001001",
				"011010011010",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"010010011000",
				"010010011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010001111000",
				"010001110111",
				"010001100110",
				"010001010101",
				"001101000101",
				"010001100111",
				"010110001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010001110111",
				"010110001000",
				"110011101110",
				"111011111111",
				"110111111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011101111",
				"111111111111",
				"111011101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110011101110",
				"110011111110",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011101111",
				"101111101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101110",
				"101011001100",
				"101111011101",
				"101011011101",
				"101011011101",
				"101011001100",
				"101011001100",
				"101111001101",
				"110011001101",
				"110111011101",
				"111011011110",
				"110111011101",
				"110111011101",
				"111011011110",
				"110111001101",
				"110010111100",
				"110111011110",
				"110011001101",
				"110011011101",
				"110111011110",
				"110011011110",
				"101111001101",
				"101111011101",
				"101111011110",
				"101111001101",
				"101111001101",
				"110011001101",
				"101010111100",
				"101010111100",
				"101011001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011110",
				"011111001101",
				"011010111101",
				"011011001101",
				"011111011110",
				"100011011111",
				"100011011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011011110",
				"110111011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011011101",
				"110111011101",
				"110111011101",
				"110011011100",
				"110011001100",
				"110011011100",
				"101111011100",
				"101011001100",
				"100110111011",
				"100110111100",
				"100111001100",
				"100111001100",
				"100011001101",
				"100111001101",
				"100011001101",
				"100011001100",
				"011110111100",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011011100",
				"011111011101",
				"011111011101",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110101100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011011001100",
				"010111001100",
				"010111001101",
				"011011011101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"100010111101",
				"011110111100",
				"011110101100",
				"011010101100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011011011101",
				"011011011101",
				"011011011110",
				"011111001110",
				"011111001101",
				"011010111101",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110001001",
				"010001100110",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110011",
				"010110001000",
				"011010101010",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"100111001110",
				"100010111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100111011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011011110",
				"011011011110",
				"011011011110",
				"011011001101",
				"100011001101",
				"100111001110",
				"101011001101",
				"101010111100",
				"100010011010",
				"011110001001",
				"100110111100",
				"101011001101",
				"101011011101",
				"100011011101",
				"011111011101",
				"011111011101",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100110111100",
				"100111001101",
				"101011001101",
				"100110111101",
				"101111011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100011011101",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010101010",
				"011110101011",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011001",
				"011010101010",
				"011110101011",
				"011110111011",
				"100010111011",
				"100010101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001100111",
				"010001010110",
				"001101010101",
				"010001100110",
				"010001110111",
				"010110001000",
				"011010001001",
				"010110001000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101100111",
				"010001110111",
				"010001110111",
				"001101110110",
				"010110001000",
				"101011011101",
				"110011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111111111111",
				"111011101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"101111101110",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101110",
				"110111101110",
				"110111011110",
				"101111011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011001101",
				"110010111100",
				"101110011010",
				"101010011001",
				"101010011001",
				"101110011010",
				"101110011010",
				"101010011001",
				"100110001000",
				"100110001001",
				"101010001001",
				"101010001001",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101011",
				"101110101011",
				"101110101100",
				"100110011010",
				"101010101011",
				"101110111101",
				"101111001101",
				"101111001110",
				"101011001101",
				"101011001101",
				"101011001110",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100011001101",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001100",
				"110011011101",
				"110011011100",
				"110011011101",
				"110111011101",
				"110111011101",
				"110011011100",
				"101111001100",
				"101111001100",
				"101111001100",
				"100110111011",
				"100110111011",
				"100111001100",
				"101011011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100011001101",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011110111100",
				"100011001100",
				"100011001101",
				"100010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011111001100",
				"011111001101",
				"011011001101",
				"011011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011110111100",
				"011110101100",
				"011010101100",
				"011110111100",
				"011111001101",
				"011011001100",
				"011010111100",
				"011011001100",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110001001",
				"010001100110",
				"000100100011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101010101",
				"010110001000",
				"011010101010",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111101",
				"100010111100",
				"100010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111001101",
				"100011001101",
				"100111001110",
				"101011001101",
				"100110101100",
				"011110011010",
				"011010001001",
				"011110101011",
				"100010111100",
				"100111001101",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111011101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"101011011101",
				"101011001101",
				"100110111100",
				"100110111100",
				"100110111100",
				"101011001101",
				"101011001101",
				"100111001101",
				"101011011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010011010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"001101110111",
				"001101110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010110001000",
				"011110101010",
				"101111011101",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111111111111",
				"111011101111",
				"111011101110",
				"111011101111",
				"110111101110",
				"110111101110",
				"110111101110",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101111",
				"101111011110",
				"110011101110",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111101110",
				"110011011101",
				"110111011110",
				"111011101110",
				"110111101110",
				"110011011101",
				"101111001100",
				"101010111011",
				"101110111011",
				"101110101011",
				"101010011010",
				"100110001000",
				"100001110111",
				"100001100110",
				"011101010101",
				"010100110100",
				"001100010010",
				"001100010010",
				"011001000100",
				"100101110111",
				"100001110111",
				"010101000100",
				"010000110100",
				"011001010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101111000",
				"011101111000",
				"011001100111",
				"011101111000",
				"100110011010",
				"101010101011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101110111101",
				"101111001101",
				"101111001110",
				"101111001110",
				"101111001101",
				"101011001101",
				"101111011110",
				"100111011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011011101",
				"100111011101",
				"100111011110",
				"101011011110",
				"100111011110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011001100",
				"110011011100",
				"110011011100",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011011100",
				"101111001100",
				"101111001100",
				"101011001100",
				"100110111011",
				"100110111011",
				"101011001101",
				"101011011101",
				"101011011101",
				"100111001101",
				"100111001101",
				"100011001100",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011011001100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111011101",
				"011011011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011010111100",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011011001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110001001",
				"010001100110",
				"000100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001000100",
				"010001110111",
				"010110011010",
				"011010101011",
				"011110111100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011110111100",
				"100010111101",
				"100010111100",
				"100010101100",
				"100010101011",
				"100010011011",
				"100010101011",
				"100010101100",
				"100010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011001110",
				"011111001110",
				"100111001110",
				"100111001110",
				"100010111100",
				"011110011011",
				"011110011010",
				"011110101011",
				"011110111011",
				"100011001101",
				"100011011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011111",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111001101",
				"101010111100",
				"100110101011",
				"100110101011",
				"100110101011",
				"101011001100",
				"101011001101",
				"100111001101",
				"100111011101",
				"100011001101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011001110",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011011101",
				"100111011101",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"100111001101",
				"100010111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011111001100",
				"011010111011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111100",
				"011110101011",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111010",
				"011010101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010010011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"011010101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"001101110111",
				"010010001000",
				"010001110111",
				"001101110110",
				"001101100110",
				"011110101010",
				"110011101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011101111",
				"111011101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"111011101111",
				"111011111111",
				"111011101111",
				"110111101111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101110",
				"101111011110",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110011001101",
				"101010101010",
				"101010101010",
				"101010101010",
				"100010011001",
				"100010011001",
				"100010001001",
				"011110001000",
				"011101100111",
				"011101010110",
				"011001010110",
				"011001000101",
				"101010011001",
				"101010011001",
				"011001100101",
				"010000110011",
				"010000110011",
				"010001000100",
				"011001010101",
				"101010101010",
				"101110101010",
				"011101110111",
				"011001100110",
				"100010001000",
				"100110101010",
				"100110011010",
				"100110101010",
				"100110111011",
				"100110101010",
				"011110011001",
				"011110001000",
				"100010011001",
				"100010011001",
				"011101111001",
				"011110001001",
				"100010001001",
				"101010101011",
				"101010101100",
				"101110111100",
				"101110111100",
				"101010111100",
				"101010111011",
				"101010111100",
				"101011001101",
				"101111011110",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"100111011101",
				"100111011101",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101111001101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011011100",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100111001100",
				"101011001100",
				"101011001101",
				"100111001100",
				"100111001101",
				"100111011101",
				"011110111100",
				"011010101011",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001011",
				"011111001100",
				"011110111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011011001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001100",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110101011",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110001001",
				"010001100111",
				"000100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100110100",
				"010001100111",
				"011010011010",
				"011010101011",
				"011110111100",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011011011101",
				"011111001101",
				"100011001101",
				"100110111101",
				"100010011011",
				"100010011011",
				"100010001010",
				"100110101100",
				"100010111100",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011001110",
				"100111001110",
				"100111001110",
				"100010111101",
				"100010111100",
				"100010111101",
				"100111011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111001110",
				"101011011110",
				"101011011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011001110",
				"100110111101",
				"100110101100",
				"100010001001",
				"100010001001",
				"100010011010",
				"101010111100",
				"101011001101",
				"100111011101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011110111100",
				"100011001101",
				"100111001101",
				"100111001101",
				"100110111101",
				"100110101100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011110101010",
				"011110111011",
				"011010111011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010101010",
				"010010011010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"001101111000",
				"001110001000",
				"010010001001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010010001000",
				"010001110111",
				"011010011001",
				"100111001100",
				"110011111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101110",
				"111011101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011101110",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101110",
				"110011011101",
				"101111001100",
				"101010101011",
				"100110011001",
				"100110011001",
				"100010011001",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110101011",
				"101110101011",
				"101010011010",
				"100110011001",
				"101110111011",
				"101010111011",
				"100110101010",
				"100110011010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101111011101",
				"110011011101",
				"110011101110",
				"101111011110",
				"101111011101",
				"101111101101",
				"101011011101",
				"101011011100",
				"101111011101",
				"101010111100",
				"100010011010",
				"100010011010",
				"100010001001",
				"011101111001",
				"100010001001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100110111011",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011101",
				"100111011101",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011011100",
				"110011011100",
				"101111011100",
				"101111001100",
				"101011001011",
				"100110111011",
				"100110111011",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001100",
				"101011011101",
				"011110111011",
				"011010111011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011111001100",
				"011110111011",
				"011010111011",
				"011010101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111011101",
				"100011011101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"011110101011",
				"011110101011",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110101100",
				"011010101011",
				"011110101100",
				"011110101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110001001",
				"010001110111",
				"000100110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000101000100",
				"010001100111",
				"011010011010",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111011110",
				"011011011110",
				"011011011101",
				"100011011110",
				"100111001110",
				"100110111101",
				"100110101100",
				"100110011011",
				"100010011011",
				"101010111101",
				"100111001101",
				"100011001101",
				"100011011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011001110",
				"100010111101",
				"100010111101",
				"100111001110",
				"100111011111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011011111",
				"100111011110",
				"100111001110",
				"100011001101",
				"100010111101",
				"100010111101",
				"100110111101",
				"100110111101",
				"100110111101",
				"100110111100",
				"100010101011",
				"100010011010",
				"011110001001",
				"011101111000",
				"011101111001",
				"100010001010",
				"100110101011",
				"100111001100",
				"100111011101",
				"100011011101",
				"011111001101",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011010111101",
				"011010111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100110101100",
				"100010011011",
				"011110011010",
				"011110101011",
				"100010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011001111000",
				"010101100111",
				"010101100111",
				"011001111000",
				"011110011010",
				"011110101011",
				"011110111011",
				"011010111011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010110101001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010101010",
				"010010101010",
				"010010101010",
				"010010101010",
				"010110101010",
				"010010011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001000",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110101010",
				"010110011001",
				"010010011001",
				"010010011000",
				"010010001000",
				"010010001000",
				"010010000111",
				"010001110111",
				"010010001000",
				"010110001001",
				"010010001000",
				"010010001000",
				"001101111000",
				"001101111000",
				"001101111000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010001110111",
				"010110001000",
				"010001110111",
				"010001111000",
				"011110101010",
				"101011011101",
				"101111101110",
				"110011111111",
				"110011101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"111011101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110111101110",
				"110111101110",
				"101111001101",
				"101110111100",
				"100110011010",
				"100110011010",
				"101010101010",
				"101110111011",
				"110111011101",
				"110111101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111011110",
				"101111001101",
				"100110111100",
				"100111001100",
				"101111101110",
				"101111101110",
				"100111001100",
				"101011001101",
				"101111101110",
				"101111011110",
				"100111001100",
				"100111001101",
				"101011001101",
				"100111001100",
				"100011001100",
				"100111001100",
				"100111001101",
				"100011001100",
				"100011001100",
				"100011011100",
				"100111011101",
				"101011101110",
				"100111011101",
				"100111001100",
				"101011001101",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010101011",
				"100010101010",
				"011110011001",
				"011010001000",
				"011010001000",
				"100010101010",
				"100110111011",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101011011101",
				"101011011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011011101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011011100",
				"101111001100",
				"101111001011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101011001100",
				"101011001101",
				"101011001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001100",
				"100111001100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"100011001100",
				"011110111011",
				"011010101011",
				"011010101010",
				"011010111011",
				"011011001011",
				"011011001011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111011101",
				"100011011101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011011101",
				"011111011101",
				"011111011101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110101100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011110101100",
				"011110101011",
				"011110101100",
				"011110101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011001",
				"010001110111",
				"001000110100",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100110011",
				"001101100111",
				"010110011001",
				"011010101011",
				"011110111100",
				"011110111101",
				"011111001101",
				"011010111101",
				"011110111101",
				"011111001101",
				"100011001110",
				"100011001101",
				"100011001110",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011011110",
				"011011011110",
				"011011011110",
				"100011011110",
				"100111001110",
				"100110111101",
				"100110101100",
				"100110011100",
				"100110101100",
				"101011001101",
				"100111001101",
				"100011001101",
				"011111011101",
				"011111011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"100111001110",
				"100111011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111011111",
				"100011011111",
				"100011011111",
				"100111011111",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111101",
				"100010111100",
				"100010101100",
				"100010011011",
				"100010001010",
				"100010001010",
				"100010001001",
				"100110011010",
				"100110111100",
				"101011001101",
				"100111001101",
				"011111001100",
				"011011001100",
				"011011011101",
				"011011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100110111101",
				"101010111101",
				"101010101100",
				"100110101011",
				"100110101011",
				"100110111100",
				"100111001101",
				"100011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011110101011",
				"011110101010",
				"011110011010",
				"100010011010",
				"011101111001",
				"010101100111",
				"011110001001",
				"100010101011",
				"100010111100",
				"100010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110111010",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010010101010",
				"010010011010",
				"010010011001",
				"010110011010",
				"010110011001",
				"010110001001",
				"010101111000",
				"010001110111",
				"010001100110",
				"001101100110",
				"010001100111",
				"010001111000",
				"010110001001",
				"011010011001",
				"010110011001",
				"010010011001",
				"010010001000",
				"001110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010011001",
				"010010001001",
				"001101110111",
				"001001100111",
				"001101111000",
				"010010001001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001111000",
				"010110001001",
				"100011001100",
				"100111011101",
				"101111101110",
				"101111011110",
				"110111101111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101110",
				"110011011101",
				"101111001100",
				"101010101011",
				"100010011010",
				"100110101010",
				"101010101011",
				"110011001101",
				"110111101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011101110",
				"101111011110",
				"101111011101",
				"100111001101",
				"101011011110",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111011110",
				"100111001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011100",
				"100011011101",
				"100111011101",
				"100111011101",
				"100011001100",
				"100011001100",
				"100111001101",
				"100010111100",
				"100010111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011001101",
				"100010111011",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100110111011",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101011011101",
				"100111011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101111011101",
				"101111011101",
				"101111001100",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011011100",
				"101111001100",
				"101011001011",
				"100110111011",
				"100110111011",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001101",
				"101011001100",
				"100111001100",
				"100111001100",
				"101011011100",
				"100111001100",
				"100010111011",
				"011010101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011111001011",
				"011110111011",
				"011110111011",
				"100011001100",
				"100011001100",
				"011110111011",
				"011010101011",
				"011110111011",
				"011111001100",
				"011011001011",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001100",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011011101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011111001101",
				"100011011101",
				"100011001101",
				"011110111100",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011011101",
				"011011011101",
				"011011001100",
				"011011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011110",
				"011111011101",
				"011011001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011001",
				"010001110111",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100110011",
				"010001100110",
				"011010011001",
				"011110101011",
				"011110111100",
				"011111001101",
				"011010111101",
				"011011001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011011011110",
				"011111011110",
				"100011011110",
				"100111011110",
				"100111001110",
				"100110111101",
				"100010101100",
				"100010101100",
				"100111001101",
				"100011001101",
				"100011011110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011011110",
				"100011101110",
				"100011011110",
				"100011011110",
				"100111011111",
				"100111011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100111001110",
				"100111001110",
				"100111011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011011110",
				"100011001101",
				"100010111100",
				"100110111101",
				"100110101100",
				"100110011011",
				"101010101100",
				"101010111101",
				"101011001110",
				"100111011110",
				"100011001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011011101",
				"011011011101",
				"011111011101",
				"011111001101",
				"011110111100",
				"100010111100",
				"100110101100",
				"101110111101",
				"101010101100",
				"101010111101",
				"101111011110",
				"101011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"010111001100",
				"010111001011",
				"010111001100",
				"010111001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110101011",
				"011110011010",
				"100010011010",
				"100010011010",
				"011110001001",
				"011001111000",
				"100010011010",
				"100110111100",
				"100110111100",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010111011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"011010011010",
				"010110001000",
				"010101111000",
				"001101010110",
				"001101010101",
				"010101111000",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010010001001",
				"010010011000",
				"010010001000",
				"010010011000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"001101111000",
				"001101110111",
				"001101100111",
				"010001111000",
				"010110001001",
				"010110001001",
				"010101111000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010110011001",
				"010110011001",
				"011110111011",
				"100111001101",
				"101011001101",
				"110011011110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101111",
				"111011101111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111101110",
				"101111001101",
				"101010101011",
				"100110101011",
				"101010111011",
				"101111001100",
				"110011011101",
				"110011011110",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111101110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011011110",
				"101011011110",
				"100111011101",
				"100111011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100010111100",
				"100010111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011101",
				"100111011101",
				"100011001101",
				"100011001100",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100110111100",
				"100111001100",
				"100111001101",
				"101011001100",
				"101011001100",
				"101010111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"101010111011",
				"101111001100",
				"110011011101",
				"101111001101",
				"101111011101",
				"101111011110",
				"101111011110",
				"100111011101",
				"100111011101",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011011101",
				"101111011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011011101",
				"110011011100",
				"101111001100",
				"101011001011",
				"101011001011",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011011101",
				"101011001101",
				"100111001100",
				"100110111100",
				"100111001100",
				"101011011101",
				"101011001100",
				"100110111011",
				"011110101010",
				"011010101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"100011001100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011010101010",
				"011010111011",
				"011110111011",
				"011111001011",
				"011010111011",
				"011011001011",
				"011011001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011111001100",
				"011111001101",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001101",
				"100011001101",
				"100011011101",
				"011110111100",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011011101",
				"011011011101",
				"011011011101",
				"011011011101",
				"011011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100111001101",
				"100010111101",
				"011110111100",
				"011010101011",
				"011010111011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011011001101",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"010001111000",
				"001101010101",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101010101",
				"010110001001",
				"011110101011",
				"011110111100",
				"011111001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011111",
				"100111011110",
				"100111001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100111001110",
				"100111001110",
				"100111001101",
				"100110111101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101110",
				"100011011110",
				"100011101110",
				"100011101110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100011011110",
				"100111011111",
				"100111011111",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111001110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011111",
				"011111011111",
				"011111101111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111001101",
				"100011001101",
				"101011001101",
				"101010111100",
				"101010101100",
				"101110111101",
				"101011011110",
				"100111001110",
				"100011001110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011011101",
				"011011001101",
				"011111001100",
				"011110111100",
				"100010111100",
				"100110111101",
				"101010111101",
				"100110101100",
				"100110101100",
				"101011001101",
				"100111001110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011011100",
				"010111011100",
				"010111011100",
				"010111001100",
				"010111001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110011010",
				"100010101011",
				"100010011010",
				"011001111000",
				"010001010110",
				"011010001001",
				"100010101011",
				"100111001100",
				"100011001100",
				"011110111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010010101011",
				"010010101011",
				"010110111011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110011001",
				"011010001000",
				"011010001000",
				"010101100111",
				"010001100111",
				"011110001001",
				"100010101011",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"001101111000",
				"010001111000",
				"010001100111",
				"010001101000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010110001000",
				"010110001001",
				"010010001001",
				"001110001000",
				"010110001001",
				"100011001100",
				"101111101111",
				"110011101110",
				"110111101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"110011011101",
				"101010111011",
				"100110101011",
				"101010111100",
				"110011011101",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101111",
				"101011101110",
				"100111011110",
				"100111011101",
				"100111011110",
				"101011011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001110",
				"100111001110",
				"100011001101",
				"100010111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100110111100",
				"100110101011",
				"101011001100",
				"110011011101",
				"101111001101",
				"101010111011",
				"100110101010",
				"101010101011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011011101",
				"101111011101",
				"101011001101",
				"101011011101",
				"101011011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111011101",
				"101011011101",
				"101011011101",
				"101111011100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001011",
				"101011001011",
				"101111001100",
				"101111011100",
				"101111011100",
				"101111011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"100111001100",
				"101011001100",
				"101011011101",
				"101011001100",
				"100110111011",
				"011110101010",
				"011010101010",
				"011010111010",
				"011010111011",
				"011110111011",
				"011111001011",
				"011111001011",
				"011111001100",
				"011111001100",
				"100011001100",
				"011110111011",
				"011110111011",
				"011010101010",
				"011010101010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"011110101011",
				"011010101011",
				"011010111011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011010101011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011011001100",
				"011111011100",
				"011111011101",
				"011011011101",
				"011011011101",
				"011011001101",
				"011011001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"011110111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011010101101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110001000",
				"001101010110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001000100",
				"010110001000",
				"011110101011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111011111",
				"101011011111",
				"100111001110",
				"100011001101",
				"100010111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"100011001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011101110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011011111",
				"100111001110",
				"100010111101",
				"100011001101",
				"100111011111",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101110",
				"011111011110",
				"011111011110",
				"011111001101",
				"100011001101",
				"101011001110",
				"101010111101",
				"101110111101",
				"110011001110",
				"101011011111",
				"100011011110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111101101",
				"011111101110",
				"011111101110",
				"011111011110",
				"011011011110",
				"011011011101",
				"011011001101",
				"011011001100",
				"011110111100",
				"100010111100",
				"100110111100",
				"100110111101",
				"100010011011",
				"100010011011",
				"100110111101",
				"100111001110",
				"100111011110",
				"100111101110",
				"100011011110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011011011101",
				"011011011100",
				"011011011100",
				"011011011100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010011010",
				"011110011010",
				"100010011010",
				"011110001001",
				"010101101000",
				"010001010111",
				"010101111000",
				"011010001001",
				"011110101011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010010101010",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"011010001001",
				"011110001001",
				"010101111000",
				"010001100111",
				"011010001001",
				"100010101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010101111000",
				"010001111000",
				"010001101000",
				"010001100111",
				"010001100111",
				"010101111000",
				"011010001001",
				"011010011001",
				"010010001000",
				"001101111000",
				"001101110111",
				"011110101011",
				"110011111111",
				"110011101111",
				"101111001101",
				"110111101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"101110111100",
				"101111001100",
				"101111001101",
				"110011011110",
				"110111101111",
				"111011111111",
				"110111101111",
				"110011101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101110",
				"100111101110",
				"101011101111",
				"101011111111",
				"101011101111",
				"101011101110",
				"100111011101",
				"100111011101",
				"101011011110",
				"100111011101",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100011001100",
				"100111001100",
				"100111001101",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001101",
				"101011011110",
				"100111001101",
				"100010111101",
				"100010111100",
				"100010111101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011111001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"100110101011",
				"100110111011",
				"101010111100",
				"101011001100",
				"101111001101",
				"101111001101",
				"101110111100",
				"100110101010",
				"101010101010",
				"101110111100",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101011011101",
				"101011011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011101",
				"100111011101",
				"100011001101",
				"100111001100",
				"100111001101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101111001100",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001011",
				"101011001100",
				"101111001100",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100110111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011111001011",
				"011111001011",
				"011110111011",
				"011110111011",
				"100011001100",
				"100011001100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011111011101",
				"011111011101",
				"011111011101",
				"011011011101",
				"011011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111011101",
				"100011001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101100",
				"011010111100",
				"011110111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010101010",
				"010110001001",
				"010001100110",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"001101100110",
				"011010011010",
				"011110111011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"100011001110",
				"100111011110",
				"100111011111",
				"100111001110",
				"100010111101",
				"100010111101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001101",
				"100011001110",
				"100011011110",
				"100111011110",
				"100111011111",
				"100011011111",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100111011111",
				"101011101111",
				"101011011111",
				"100110111101",
				"100010101100",
				"100010111101",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101110",
				"011111011110",
				"011111011110",
				"100011001101",
				"100111001101",
				"101011001101",
				"101010111100",
				"101010101100",
				"101010111101",
				"101011011111",
				"100011011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101110",
				"011111101110",
				"011111101110",
				"011111101110",
				"011111101110",
				"011111101101",
				"011111101110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111001100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100110111101",
				"100010101100",
				"100010111100",
				"100111001110",
				"100111011110",
				"100111011110",
				"100011101110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011011001100",
				"011011001100",
				"011111011100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010011010",
				"011110011010",
				"011110001010",
				"011110001001",
				"011110011010",
				"011110101011",
				"011110101011",
				"011010101011",
				"011110111011",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010001001",
				"011010001001",
				"010101100111",
				"001101010110",
				"010101100111",
				"011010001001",
				"011110011010",
				"011110101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010001111000",
				"010101111001",
				"011001111001",
				"010101111000",
				"010101111000",
				"011010011001",
				"011110011010",
				"010110011001",
				"010010001000",
				"010010001000",
				"001101111000",
				"010110011001",
				"101011011101",
				"110011101111",
				"101011001101",
				"101011001101",
				"110111111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110111101110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110111011110",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101111",
				"101111101110",
				"101011101110",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101011101110",
				"101011011110",
				"101011011101",
				"101011101110",
				"101011011101",
				"101011011101",
				"100111011101",
				"100111011100",
				"100111011101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100111001100",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100110111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011111001101",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"100110111011",
				"100110111100",
				"100110111100",
				"101010111100",
				"101011001100",
				"101111001100",
				"101111001100",
				"100110101010",
				"101010101010",
				"101010111011",
				"110011011100",
				"110011011101",
				"101111011101",
				"101011001101",
				"101011001101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101111001100",
				"101111011101",
				"101111011101",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101111011100",
				"101111011101",
				"101011001100",
				"100111001100",
				"100111001011",
				"100111001100",
				"100111001100",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111011",
				"100010111011",
				"100011001100",
				"011111001011",
				"011111001011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"100011001100",
				"100011001100",
				"100111011101",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011111001100",
				"100011001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001101",
				"011110111101",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011011011101",
				"011111011110",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011010111101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110001001",
				"010001100110",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001001000100",
				"010110001000",
				"011110101011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"100111011110",
				"100111001110",
				"100011001110",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100111011110",
				"101011011111",
				"101011001110",
				"100110111101",
				"100110111101",
				"100111001110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111011110",
				"100011011111",
				"100011001110",
				"100110111101",
				"100110111101",
				"101010111101",
				"100110101100",
				"100110101100",
				"100110111101",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"011111101110",
				"011111101110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011110111100",
				"100010111100",
				"100010111100",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"010110111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100110111100",
				"101011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"011010001001",
				"011010011010",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"001110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"011010001001",
				"011110011010",
				"010110011001",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001110111",
				"011010101010",
				"101011011101",
				"101111011110",
				"101011001101",
				"101111011101",
				"110011101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101110",
				"110011011110",
				"110011011110",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110011111111",
				"110111111111",
				"110011111111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011101101",
				"101011011101",
				"101011011101",
				"100111011101",
				"100111011100",
				"100111011100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111011100",
				"100111011100",
				"100111011101",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011110111100",
				"011110111100",
				"100010111011",
				"100110111100",
				"100111001100",
				"100110111100",
				"100010101011",
				"100010101011",
				"101010111100",
				"101111011101",
				"101010111011",
				"101010101010",
				"100110101010",
				"101110111011",
				"110011001100",
				"110011001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001101",
				"101011011101",
				"101011001100",
				"101011001101",
				"101111011101",
				"101111011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001011",
				"101111001100",
				"101111011100",
				"101111011100",
				"101011001100",
				"100110111011",
				"100010111011",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100010111011",
				"011110111011",
				"011010111010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100011001100",
				"100111001101",
				"100111001100",
				"100010111011",
				"011110101010",
				"011110111010",
				"011010111011",
				"011010111010",
				"011010101010",
				"011010111011",
				"011110111011",
				"011110111011",
				"011111001100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011111001100",
				"011111001100",
				"100011011101",
				"100111011101",
				"100011011101",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100111011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"100011001101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011111001101",
				"011110111101",
				"011010111101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011011001101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110111011",
				"011010101011",
				"010110011010",
				"010110001000",
				"001101100110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101010110",
				"011010011010",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111011101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011011110",
				"100011001110",
				"101011001110",
				"101011001110",
				"101010111101",
				"101111001110",
				"101111011111",
				"100111011110",
				"100011011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011001101",
				"100110111101",
				"100110111101",
				"101010111101",
				"101011001101",
				"101011001110",
				"101011011110",
				"100111011110",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100011011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"100011001101",
				"100111001101",
				"100111001110",
				"100111001110",
				"101011011111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"100011001101",
				"100011011101",
				"100111011110",
				"100111011110",
				"100011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011110101011",
				"100010101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010001101000",
				"010001100111",
				"010101101000",
				"010101111000",
				"010101111000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"001101110111",
				"010001111000",
				"011110101010",
				"101011011101",
				"101011011101",
				"101111011110",
				"101111011101",
				"110111101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101110",
				"101111011110",
				"101111011110",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011011101",
				"100111011101",
				"100111001100",
				"101011011101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111011100",
				"100111011100",
				"100111001100",
				"100111001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111100",
				"100111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100011001100",
				"011110111100",
				"011110111011",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100110111011",
				"101010111011",
				"110011011101",
				"101111001011",
				"101010101010",
				"100110101001",
				"101010101011",
				"110011001100",
				"110011011101",
				"101111011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101111011101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001011",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001100",
				"101011001011",
				"100110111011",
				"100010111011",
				"100011001100",
				"100111001100",
				"101011001101",
				"100111001100",
				"100010111011",
				"011110101010",
				"011010101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"100010111100",
				"100111001100",
				"100111001100",
				"100010111011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011111001011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011111001100",
				"011111001100",
				"100011011101",
				"100111011101",
				"100111011101",
				"100011001101",
				"011111001100",
				"011110111100",
				"011111001100",
				"100011001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011101",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100010111100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101100",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010101010",
				"010110001000",
				"001101010110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110100",
				"010001111000",
				"011110101011",
				"011110111100",
				"011111001100",
				"100011011101",
				"011111011101",
				"011111001100",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100111011110",
				"100111011111",
				"100111011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111101111",
				"011111011111",
				"100011011111",
				"100011001110",
				"100111001110",
				"101010111110",
				"101110111101",
				"110011001110",
				"110011011111",
				"101011011110",
				"100111101110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011111111",
				"100011111111",
				"011111111111",
				"011111101111",
				"011111101111",
				"100011011110",
				"100011001110",
				"100011001101",
				"100110111101",
				"101011001110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101011101111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100011101110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100111001110",
				"101011011110",
				"101011011111",
				"101111101111",
				"101011011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"011111011101",
				"011111011110",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100111011110",
				"100111011101",
				"100111011110",
				"100111011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"100011001110",
				"100011001110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011010101010",
				"011110101011",
				"011110101011",
				"100010111100",
				"100010111100",
				"011110101011",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010001111000",
				"010101111000",
				"011010001001",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010001111000",
				"001101110111",
				"010010001000",
				"011110101011",
				"101011011101",
				"110011101110",
				"110011101110",
				"110111101111",
				"111011111111",
				"111011101111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011011101",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"101011001101",
				"100111001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100011001011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"101011001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"100010111100",
				"100011001101",
				"100011001100",
				"100010111100",
				"100010111011",
				"100110111011",
				"101010111011",
				"101111011100",
				"110011011100",
				"101111001011",
				"101010101010",
				"101010101010",
				"101110111011",
				"110011001100",
				"110011011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"101011001100",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001011",
				"101111001011",
				"101111001011",
				"101111001011",
				"101011001011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100111001100",
				"101011001101",
				"101011001100",
				"100110111100",
				"011110111011",
				"011010101010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100111001100",
				"100110111100",
				"100010111011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011110111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001011",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011011101",
				"100011001100",
				"011110111011",
				"011010101011",
				"011010101010",
				"011110111011",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001011",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011011101",
				"100011011101",
				"100011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"100111011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100010111101",
				"100010111100",
				"100010101100",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011011001110",
				"011011011110",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011010111011",
				"011010101010",
				"010001110111",
				"001001000101",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100011",
				"001101010110",
				"010110001010",
				"011110111100",
				"100011001101",
				"011111001101",
				"100011011101",
				"100011011101",
				"011111001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111011110",
				"100011001110",
				"100011011110",
				"100111011111",
				"100111101111",
				"100111011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"100011011111",
				"100011001110",
				"101011001110",
				"101011001110",
				"101010101101",
				"101010111101",
				"101111011111",
				"101111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"011111111111",
				"011111101111",
				"011111101110",
				"100011011110",
				"100011011110",
				"100111001110",
				"100111011110",
				"101011011111",
				"101011101111",
				"101111111111",
				"101011111111",
				"100111101111",
				"101011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111011111",
				"100111011110",
				"100111001110",
				"100111001110",
				"101011011110",
				"101011011111",
				"101011011111",
				"101011101111",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011101110",
				"011111101110",
				"011111101110",
				"100011101111",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110111100",
				"100111011110",
				"100111011111",
				"100111001101",
				"100011001101",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"011110101010",
				"011010011010",
				"011110101011",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011010",
				"010110101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010110001001",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"001101110111",
				"010110011001",
				"100111001100",
				"101111101110",
				"110011101110",
				"110111111111",
				"111011111111",
				"110111011110",
				"110111101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"101111111111",
				"101111101111",
				"101111101110",
				"101111101110",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111111111",
				"110111101111",
				"110111101110",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011001101",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011001100",
				"100111001100",
				"101011001101",
				"100111001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001100",
				"100110111100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"100010111100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111011",
				"100010111100",
				"100110111100",
				"100110111011",
				"101010111011",
				"101111001100",
				"110011011100",
				"110011001100",
				"101010101010",
				"100110011001",
				"101010101010",
				"101111001100",
				"101111001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"101111001100",
				"101111001011",
				"101011001011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100111001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"011110111011",
				"011010111010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"100010111011",
				"100111001100",
				"100110111011",
				"100010111011",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011111001011",
				"011111001100",
				"011110111011",
				"011110111011",
				"011111001100",
				"100011001101",
				"100011001100",
				"011110111011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110111010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011111001011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001011",
				"011111001100",
				"100011011101",
				"100111011101",
				"100011001101",
				"100010111100",
				"011110111011",
				"011010111011",
				"011110111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"100011011101",
				"100011011101",
				"100111011110",
				"101011011110",
				"100111011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111001101",
				"011010111101",
				"011010111100",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111101",
				"100010111101",
				"100011001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011010111011",
				"010110011010",
				"001101100111",
				"000100110100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001101010101",
				"010110001000",
				"011010101011",
				"011010111100",
				"100011001101",
				"100011011110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001110",
				"011111011110",
				"011111011110",
				"011011011110",
				"011111011110",
				"100011011110",
				"100111011111",
				"100111011111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"011111011110",
				"011111011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111001110",
				"100111001110",
				"100010111101",
				"100011001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100111011110",
				"100111001110",
				"100111001110",
				"101011001110",
				"101011011111",
				"101011011110",
				"100111011111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101110",
				"100011111111",
				"100011111111",
				"100011101110",
				"100011101110",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"101011011111",
				"101011011111",
				"101011001110",
				"100111001101",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010111101",
				"101011011110",
				"101011101111",
				"100111101111",
				"100011011110",
				"100011011110",
				"100011101111",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110101011",
				"011110011011",
				"011110011010",
				"011110001010",
				"011110001001",
				"011010011010",
				"100010111101",
				"100011001101",
				"100111011110",
				"100011001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010101100",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011110101010",
				"011110011010",
				"011110001001",
				"011010001001",
				"011010001001",
				"011110011010",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011010011010",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001000",
				"010110011001",
				"010010001000",
				"001101110111",
				"010010001000",
				"011110101010",
				"101111101110",
				"110011101111",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"111011101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"101111101110",
				"101111011110",
				"110011101111",
				"110011101111",
				"110011101110",
				"110011101110",
				"110111101111",
				"110011101110",
				"110011011101",
				"110111101110",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"101111101110",
				"101111101110",
				"101111101110",
				"101111101111",
				"101011101110",
				"101011011101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011011101",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011001101",
				"100111001100",
				"100111001100",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011011101",
				"101011001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110101010",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100010111100",
				"100110111100",
				"100111001100",
				"100110111100",
				"100110111011",
				"101011001100",
				"101010111011",
				"101010111011",
				"101111001100",
				"110011011101",
				"101010111011",
				"100010011001",
				"100010011001",
				"101010111011",
				"101011001100",
				"101011001100",
				"101011001011",
				"101011001100",
				"101111001100",
				"101111001100",
				"101010111011",
				"101010111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"101111001100",
				"101010111011",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100111001100",
				"100111001100",
				"100011001011",
				"100010111011",
				"011110111011",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100111001011",
				"100111001011",
				"100111001011",
				"100010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111011",
				"011110111011",
				"011110111010",
				"011110111010",
				"011110111011",
				"011111001011",
				"011111001011",
				"011111001011",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100111001100",
				"100111001101",
				"100111001100",
				"100010111100",
				"011110111011",
				"011110111100",
				"100011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"100011011101",
				"100011011101",
				"100111011101",
				"100111011110",
				"100111011101",
				"100111001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011101",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100011001110",
				"100011001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011010111011",
				"010110011001",
				"001101100110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"010001110111",
				"010110011010",
				"011010111011",
				"011110111101",
				"011111001101",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100111011111",
				"100111011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111011111",
				"100011011111",
				"100011001110",
				"100011001110",
				"100111001111",
				"101011001111",
				"101011001110",
				"100110111101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101110",
				"011111101110",
				"011111101110",
				"011111101110",
				"011111101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011001110",
				"100111001110",
				"100111011111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101110",
				"100011011110",
				"100111101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100011111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100011001110",
				"100111001110",
				"100110111101",
				"100110111101",
				"100110101100",
				"100010011010",
				"011110001001",
				"011110011010",
				"100111001101",
				"101011101111",
				"100111101111",
				"100011011110",
				"100011101110",
				"011111011110",
				"011111101111",
				"011111101111",
				"011111011111",
				"011111011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011010101011",
				"011110011010",
				"100010011010",
				"100010001010",
				"011101111001",
				"011110001001",
				"100010011011",
				"100111001101",
				"100111011110",
				"100011011110",
				"100011001101",
				"011111001100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011001",
				"010110001001",
				"010110001000",
				"010101110111",
				"010101100111",
				"011001111000",
				"011010001001",
				"100010101011",
				"100010111100",
				"011010111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011110101011",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010001110111",
				"010001110111",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"101011001101",
				"110111111111",
				"111011111111",
				"110111101111",
				"110111011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110111101110",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110011101111",
				"101111101111",
				"101011101110",
				"101011011110",
				"101011011110",
				"101111101110",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101110",
				"101111101110",
				"101111011110",
				"101111011110",
				"101011011101",
				"100111001101",
				"101011011101",
				"101011011101",
				"101011001101",
				"101011001100",
				"101011001101",
				"101011001101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"101010111011",
				"101011001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"101011001100",
				"101111011101",
				"101111001100",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001100",
				"101111001101",
				"101111001100",
				"101111001100",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001011",
				"101010111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011010101010",
				"011010101010",
				"011110111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111010",
				"011110111010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100111001100",
				"100010111100",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011111001011",
				"100011001011",
				"100011001011",
				"100011001011",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001100",
				"100111001100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011101",
				"100111011101",
				"100111001101",
				"100011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011011001101",
				"011011001110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011011001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010011001",
				"001101010110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001000101",
				"010110001001",
				"011010101011",
				"011110111100",
				"011111001101",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100111011111",
				"100011011111",
				"100011011110",
				"011111011110",
				"011111011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100111001111",
				"101011011111",
				"101011011111",
				"101011001111",
				"100111001110",
				"100011011110",
				"100011011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011111",
				"100111101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"100010111101",
				"100010111101",
				"101011011110",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011111111",
				"011111101111",
				"011111011110",
				"011111011110",
				"100011001110",
				"100010111101",
				"100110111101",
				"100110101100",
				"100110101011",
				"100010011010",
				"101010111101",
				"101111011111",
				"101111101111",
				"101011101111",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011011001101",
				"011011001100",
				"011111001101",
				"011110101100",
				"100010101100",
				"100110101011",
				"100010001010",
				"011101111001",
				"100110011011",
				"101011001101",
				"100111011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"010110111011",
				"011010111011",
				"011010101010",
				"010110011001",
				"011010001001",
				"011010001001",
				"011001111000",
				"010101100111",
				"011110001001",
				"100110111100",
				"100111001101",
				"011110111100",
				"010110101010",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001001",
				"010110001001",
				"010101111000",
				"010001111000",
				"010001110111",
				"010010001000",
				"010110011001",
				"011010101010",
				"011110101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001110111",
				"001101110111",
				"001101110111",
				"010010001000",
				"010010001000",
				"010110001000",
				"010001110111",
				"100010101010",
				"110011011110",
				"111111111111",
				"111011111111",
				"110111101111",
				"111011101111",
				"110111101110",
				"110011011110",
				"110111101110",
				"110111101111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110011101110",
				"101111001101",
				"101111001101",
				"101111011101",
				"110011011101",
				"101111001101",
				"110011001101",
				"110111101110",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"111011111111",
				"110011101111",
				"101111101111",
				"101111101110",
				"101011011110",
				"101011011101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101111011101",
				"101111011101",
				"101111011101",
				"101011011101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101011001011",
				"101011001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001101",
				"101011001100",
				"101010111011",
				"101010111011",
				"101011001011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011011101",
				"110011001101",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"101111001100",
				"101111001100",
				"101010111011",
				"100110111011",
				"100110111011",
				"101011001011",
				"101011001100",
				"101011001011",
				"100110111011",
				"100010111011",
				"011110101010",
				"011110101010",
				"011110111010",
				"011110101010",
				"011010101010",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100010111010",
				"100010101010",
				"011110101001",
				"011110111010",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100011001011",
				"100011001011",
				"100011001011",
				"100011001011",
				"100011001100",
				"100011001100",
				"100011001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001100",
				"101011001100",
				"100110111100",
				"100010111011",
				"100010111011",
				"011111001100",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100011001100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001110",
				"011011001110",
				"011011001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001110",
				"100111001110",
				"100011001101",
				"011110111100",
				"011110101100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110001001",
				"001101010101",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"010001100110",
				"011010011010",
				"011110111100",
				"011111001101",
				"011111001101",
				"100011001110",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100111011111",
				"100111011111",
				"101011011111",
				"101111011111",
				"101011011111",
				"100111011111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011011111",
				"100011101111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111001101",
				"100110111100",
				"100010101100",
				"100110111100",
				"101011011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100011111111",
				"100011111111",
				"011111111111",
				"011111101111",
				"011111101110",
				"100011101111",
				"100011011111",
				"100011001101",
				"100110111101",
				"101010111101",
				"100110011011",
				"100110101011",
				"110011011111",
				"110011101111",
				"101011011110",
				"100111011110",
				"100011011110",
				"100011101110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011011001101",
				"011011001100",
				"011010111100",
				"011110111100",
				"011110101011",
				"100010101100",
				"100110011011",
				"011101111001",
				"100010001010",
				"101010111100",
				"101111011110",
				"100011001101",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010110111100",
				"010110111011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011110001001",
				"011110001001",
				"011001111000",
				"011101111000",
				"100110101011",
				"101010111100",
				"100010111100",
				"011110111011",
				"010110101011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010101111000",
				"010101111000",
				"010001100111",
				"001101100111",
				"010001110111",
				"010110001001",
				"011010101010",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"001101110111",
				"001001100110",
				"001001100110",
				"010001110111",
				"010110001000",
				"010110001000",
				"010101111000",
				"101010111100",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101110",
				"110111101111",
				"110111111111",
				"110111101111",
				"110111101110",
				"110011101110",
				"110111101110",
				"110011101110",
				"110011101110",
				"110111101111",
				"110111101110",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101110111100",
				"110111101111",
				"111111111111",
				"111011111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011110",
				"110011011110",
				"101111011101",
				"101111001101",
				"101111001101",
				"101011011101",
				"101011001101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101011001100",
				"101011001100",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"100110111100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101011001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111100",
				"101110111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"100010101011",
				"011110011010",
				"100010101010",
				"100010101011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"101011001100",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101010111011",
				"101010111011",
				"101111001100",
				"101111001100",
				"101010111011",
				"101110111011",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001011",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101111001100",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"101011001011",
				"101011001100",
				"101010111011",
				"100110111011",
				"100010101010",
				"011110101010",
				"011110101010",
				"100010111011",
				"011110111011",
				"011110101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111010",
				"100010101010",
				"011110011001",
				"011110101010",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111011",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111011",
				"100010111011",
				"100010101010",
				"100010101010",
				"100010111011",
				"100010111011",
				"100011001011",
				"100011001011",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"100110111011",
				"100010101010",
				"011110111011",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"100011001101",
				"100011011101",
				"100111011101",
				"100111011101",
				"100111011101",
				"100111001101",
				"101011001101",
				"101011011101",
				"100111011101",
				"100111001101",
				"100011001100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110001000",
				"001101010101",
				"000000010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001000101",
				"010110001000",
				"011110101011",
				"011110111100",
				"011111001101",
				"011111001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100111011111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111101111",
				"100111011111",
				"100011011110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100111011111",
				"100111001110",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100011111111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111001110",
				"100110111101",
				"100110101100",
				"100110101100",
				"101011001110",
				"101111011111",
				"101011101111",
				"100111101111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100011111111",
				"100011111111",
				"100011111111",
				"011111101110",
				"011111101110",
				"011111101111",
				"011111011110",
				"011111001101",
				"100010111101",
				"101010111101",
				"100110101100",
				"100110101100",
				"110011101111",
				"110011101111",
				"101011011110",
				"101011101111",
				"100111011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"011111101110",
				"011111101110",
				"011111011110",
				"011111011101",
				"011011011101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011110111100",
				"011110011011",
				"100010011011",
				"100010001010",
				"100001111001",
				"100010011010",
				"101010111101",
				"101011011110",
				"100111011101",
				"100011011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010110111100",
				"010110111011",
				"010110111011",
				"011010101011",
				"011010101010",
				"011110011001",
				"011101111001",
				"011101111000",
				"011001111000",
				"100010011010",
				"101010111101",
				"100110111100",
				"011110111011",
				"011110111100",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010110001001",
				"011010001001",
				"010101111000",
				"010001100111",
				"010101111000",
				"011010011010",
				"011110101011",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"001101111000",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100111",
				"010001100111",
				"010001100111",
				"100010011010",
				"110011011110",
				"111111111111",
				"111111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101110",
				"110111101111",
				"110111111111",
				"110111101111",
				"110011101110",
				"110011101110",
				"110011101110",
				"110011011110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110011011101",
				"101111001100",
				"101110111100",
				"101010111100",
				"101110111100",
				"110011001101",
				"111011101111",
				"111111111111",
				"111011111111",
				"111011101111",
				"110111101111",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011011101",
				"110111011110",
				"110011011110",
				"110011011101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111011101",
				"101111011101",
				"101011001100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101011001100",
				"101010111011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101010111011",
				"101010111011",
				"101011001100",
				"101010111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"101010111011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110101011",
				"100010101010",
				"100010011010",
				"100010101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"101011001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101111001100",
				"101111001100",
				"101110111011",
				"101111001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101111001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"100110111011",
				"100110111010",
				"100010101010",
				"100010101010",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"011110011001",
				"100010101010",
				"100010111010",
				"100010111011",
				"100110111011",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010111011",
				"100010111011",
				"100010111011",
				"100111001011",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"101011001101",
				"100111001100",
				"100110111100",
				"100110111100",
				"101011001100",
				"101011001100",
				"100110111011",
				"100010101010",
				"011110111011",
				"011110111011",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"100011001101",
				"011111001100",
				"100011001101",
				"100111011101",
				"100111011101",
				"100111001101",
				"101011011101",
				"101011001101",
				"101011001101",
				"101011011110",
				"100111001101",
				"100011001100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011111001100",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011110111100",
				"011110111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110101010",
				"010110001000",
				"001001000101",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100011",
				"010001100111",
				"011010011010",
				"011110111011",
				"011110111100",
				"011111001101",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011001110",
				"100011001110",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100011011110",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100111001110",
				"100111011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100111011110",
				"101011011110",
				"101011001101",
				"101010101101",
				"101110111101",
				"110011011111",
				"101111101111",
				"101011101111",
				"100011101111",
				"011111111111",
				"011111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111111111",
				"100011111111",
				"100011101111",
				"011111101110",
				"011111101110",
				"011111011110",
				"011111011110",
				"011110111101",
				"100110101101",
				"101010111101",
				"101010101100",
				"100110101011",
				"101111011110",
				"110011101111",
				"101111101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"011111101110",
				"011111011110",
				"011011011101",
				"011011011101",
				"011011011101",
				"011011001101",
				"011010111100",
				"100010111100",
				"100010101011",
				"100110011011",
				"100110011011",
				"011101111001",
				"011101111001",
				"100010101011",
				"101011001101",
				"100111101110",
				"100011101110",
				"100011011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010111001100",
				"010110111011",
				"010110101011",
				"011010101010",
				"011010011010",
				"011110001010",
				"011101111001",
				"011101111000",
				"011101111001",
				"011101111001",
				"100110101011",
				"100111001101",
				"100011001100",
				"011111001100",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010110001001",
				"011001111000",
				"011001101000",
				"011001111000",
				"011110011010",
				"011110101011",
				"011110101011",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"001101111000",
				"001101111000",
				"001101111000",
				"001101110111",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001010110",
				"010101100111",
				"100010011010",
				"110011011110",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101110",
				"110011101110",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101110",
				"110111101110",
				"110011101110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"101111001101",
				"101110111100",
				"101010111011",
				"101110111100",
				"110011001101",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011111111",
				"110111011110",
				"110011011110",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110011011110",
				"101111011101",
				"101111001101",
				"110011001101",
				"110011011101",
				"110111011110",
				"110111011110",
				"110111101110",
				"110111101110",
				"110111011101",
				"110011011101",
				"101111001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111011101",
				"101111001100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101111001100",
				"101010111011",
				"100110111010",
				"101010111011",
				"101111001100",
				"101010111100",
				"101010111011",
				"101010111100",
				"101010111011",
				"101010111100",
				"101011001100",
				"101011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101111001100",
				"110011001100",
				"101111001100",
				"101110111100",
				"101010101011",
				"100110101011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101010111100",
				"101011001100",
				"101010111011",
				"101010111011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"101111001011",
				"101111001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110101011",
				"100010101011",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100111001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101001",
				"100010101010",
				"100110111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111100",
				"101010111100",
				"101011001100",
				"101010111100",
				"100010101011",
				"011110111011",
				"011110111011",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100111001101",
				"100111001101",
				"100111001100",
				"101011001101",
				"101011001100",
				"101011001101",
				"101011001101",
				"100111001100",
				"100010111100",
				"011110111011",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110011010",
				"010001110111",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100110100",
				"010110001000",
				"011110101011",
				"011110111100",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101011101111",
				"100111011110",
				"100111011110",
				"101011101111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100111001110",
				"101011001110",
				"101010101101",
				"101010111101",
				"110011011111",
				"110011101111",
				"101011101111",
				"100011101111",
				"011111111110",
				"011111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011110111100",
				"100110101100",
				"101010101101",
				"100010101011",
				"100010101011",
				"101011001101",
				"101111101111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101110",
				"100011101110",
				"100011011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011011001101",
				"011110111100",
				"011110101100",
				"100010101011",
				"100110011011",
				"100010001010",
				"011101111001",
				"011001111001",
				"100010101011",
				"101011011110",
				"100111101110",
				"100011101110",
				"100011011110",
				"100011011101",
				"100011011101",
				"011111011101",
				"011111011101",
				"100011011101",
				"100011011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"010110111011",
				"011010101011",
				"011010011010",
				"011110011010",
				"011110001010",
				"011110001001",
				"011101111001",
				"010101010111",
				"001101010110",
				"011010001001",
				"100111001101",
				"100111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010110001001",
				"010101101000",
				"011001101000",
				"011001111001",
				"100010011010",
				"100010101011",
				"011110101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"001110001000",
				"001101111000",
				"001101110111",
				"001101110111",
				"001101100111",
				"010001100111",
				"010001100110",
				"010001010110",
				"010001010101",
				"010101110111",
				"100010101010",
				"101111011101",
				"110111111111",
				"110111111111",
				"110011101110",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101110",
				"110111101110",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001100",
				"101110111100",
				"101110111100",
				"110011001101",
				"110011011110",
				"110111101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"111011101111",
				"110111011110",
				"110011011101",
				"110111101110",
				"110011011110",
				"110011101110",
				"110011101110",
				"110011101110",
				"110011011110",
				"110011011101",
				"110011011110",
				"110111011110",
				"111011011110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"110111011110",
				"110111011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101010111011",
				"101010101011",
				"101010111011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101011001100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101111001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011011101",
				"110111011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001011",
				"101110111010",
				"101111001011",
				"101111001011",
				"101110111011",
				"110010111011",
				"101110111011",
				"101010101010",
				"101010111010",
				"100110101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100010111011",
				"100010111011",
				"100010101010",
				"100010101011",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110111011",
				"100110101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100010101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100011001100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"101010111100",
				"101010111100",
				"101011001101",
				"100111001100",
				"100010111011",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100111011110",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110011001",
				"010001100110",
				"001000110011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000101000100",
				"010110001001",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011011111",
				"100111011111",
				"100111011110",
				"100111001110",
				"100111011110",
				"100111101110",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"101011101111",
				"101011011110",
				"100011001101",
				"100011001101",
				"100111101110",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"011111101111",
				"100011101111",
				"100111101111",
				"100011001110",
				"100111001101",
				"100110111101",
				"100110101100",
				"100110101100",
				"101111001110",
				"110011101111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100011011110",
				"100011001101",
				"100010101100",
				"100110011100",
				"100110011100",
				"101011001101",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001100",
				"011110111100",
				"100010101100",
				"100110101011",
				"100010001010",
				"011110001001",
				"100010011010",
				"100110111100",
				"101011011110",
				"101111111111",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011011001100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011110101010",
				"011110011010",
				"011110001010",
				"011001111001",
				"011001101000",
				"010101101000",
				"010101111000",
				"100010101011",
				"100111001101",
				"100011001100",
				"100011001101",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110001000",
				"011001111000",
				"010101010111",
				"010101100111",
				"011010001001",
				"011110101011",
				"011110111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101010110",
				"001101010110",
				"010001100111",
				"011001111000",
				"011010001000",
				"011110011001",
				"101011001100",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"110111101110",
				"110111101110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110111011110",
				"110011101110",
				"110111111111",
				"110011011110",
				"110011001101",
				"110111101110",
				"110111101111",
				"110011011110",
				"110011011101",
				"101111001101",
				"110011011101",
				"110011011110",
				"110111101110",
				"110011011110",
				"110011011101",
				"110111011110",
				"110111011110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"110111101110",
				"110111011101",
				"110111011101",
				"110111011110",
				"110111011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101111001011",
				"101110111011",
				"101010111010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101011001011",
				"101111001011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"101110111100",
				"101010111011",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101010",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101011",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011011100",
				"110011011100",
				"101111001011",
				"101010111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110101011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100110101011",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"101010111100",
				"101111001101",
				"101011001101",
				"100110111100",
				"100010111100",
				"100010111011",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001101",
				"101011001101",
				"100111001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001110",
				"100111001110",
				"100111001101",
				"100111001101",
				"100111011110",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111011110",
				"011111011101",
				"011111011101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010101011",
				"010110011001",
				"001101010110",
				"000100100011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001010101",
				"010110011010",
				"011110111100",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100111011111",
				"100111001110",
				"100111001110",
				"100111001101",
				"100111001110",
				"101011011110",
				"101011101111",
				"101011101111",
				"100111101110",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100111011110",
				"100111001110",
				"100111001101",
				"100110111101",
				"100110101101",
				"101010111101",
				"101111001110",
				"110011101111",
				"110011111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100011101111",
				"100011101110",
				"011111011101",
				"100011001101",
				"100111001101",
				"100110101100",
				"101010101100",
				"101110111110",
				"110011111111",
				"110011111111",
				"101111111111",
				"101011101111",
				"101011101111",
				"100111101110",
				"100111101110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100010111100",
				"100110111100",
				"100110111100",
				"100110101011",
				"100010011010",
				"100010011011",
				"101010111101",
				"101111101111",
				"101111101111",
				"100111011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011011110",
				"100111011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111011",
				"011110101011",
				"011110101011",
				"100010101011",
				"011110011010",
				"011010001001",
				"011001111001",
				"011010001010",
				"100010101100",
				"100111001101",
				"100111011110",
				"100111011101",
				"011110111100",
				"011110111011",
				"011110111100",
				"100011001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110001001",
				"010110001000",
				"010110001000",
				"011001111000",
				"010001010111",
				"010001010110",
				"010101111001",
				"011110101011",
				"011110111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001010110",
				"010001100110",
				"011001111000",
				"011110001001",
				"010101110111",
				"010101110111",
				"011110101010",
				"101111101110",
				"110111111111",
				"110111101111",
				"110111011110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011101111",
				"111011111111",
				"111011101110",
				"110111101110",
				"110111101110",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011101110",
				"110011101110",
				"110011101110",
				"110111101111",
				"110111101110",
				"110011011110",
				"110011001101",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"110011011101",
				"110011011110",
				"110011011101",
				"110111011110",
				"111011101111",
				"111111111111",
				"111011101110",
				"111011101110",
				"111011101110",
				"111011101110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"100110011001",
				"100110011001",
				"101110111011",
				"110011001100",
				"101111001011",
				"101111001100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101010101011",
				"101010111011",
				"101110111100",
				"101010111100",
				"101010111011",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101111001100",
				"110011001100",
				"110011011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011011100",
				"110011011100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001011",
				"101110111011",
				"101010111010",
				"101010111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111010",
				"100110101001",
				"100010101001",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101011",
				"100110111011",
				"100110111011",
				"100010101011",
				"100010101011",
				"100110111011",
				"100110111011",
				"101010111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"101010111011",
				"101011001100",
				"101111001100",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101011001100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101111001101",
				"101111001101",
				"101011001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010111011",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011101",
				"100011011110",
				"011111011101",
				"011111001101",
				"011111011101",
				"100011011101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010101010",
				"010110001001",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101100110",
				"011010101010",
				"011111001101",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011111",
				"100111011111",
				"100111011111",
				"101011011111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111011110",
				"101011001110",
				"101011001110",
				"101011001110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"101011011111",
				"100111001101",
				"100110111101",
				"100110111101",
				"101011001110",
				"101111011111",
				"110011101111",
				"110011111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101110",
				"100011011110",
				"100011101110",
				"100111011110",
				"100111011110",
				"101011001110",
				"101111001110",
				"101111001110",
				"110011101111",
				"101111101111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100111101110",
				"100111101110",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"100111011110",
				"100111011110",
				"101011011110",
				"100111011110",
				"100111001101",
				"100111001101",
				"101010111101",
				"101110111101",
				"100110011011",
				"100010011011",
				"101111001110",
				"101111101111",
				"101011011110",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010011010",
				"011110011010",
				"011110011011",
				"100110111100",
				"100111011101",
				"100111011101",
				"100011001101",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110001001",
				"010101111000",
				"010001010111",
				"010101100111",
				"011010001001",
				"100010101011",
				"100010111100",
				"011110111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001100111",
				"001101010110",
				"001101010101",
				"001101010110",
				"010101110111",
				"011010001001",
				"011010001000",
				"010101111000",
				"010110001000",
				"100010111011",
				"110011101110",
				"111011111111",
				"110111101111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111111111111",
				"111011101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011101110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110111011110",
				"111011101110",
				"111011101110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"100110011001",
				"100110001000",
				"101110101010",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101011001011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111011",
				"101010111011",
				"101110111011",
				"101111001100",
				"101110111100",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011001",
				"100010011001",
				"100110101010",
				"101110111011",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011001100",
				"110011001011",
				"110011001011",
				"101110111011",
				"101111001011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101010111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101011",
				"100110111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"100110101010",
				"100110101001",
				"100010101001",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100110101010",
				"100010101011",
				"100010101011",
				"100110101011",
				"100110111011",
				"100010101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101111001100",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101111001100",
				"101111001101",
				"101011001100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"101010111100",
				"100110111100",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001101",
				"100111001101",
				"100111001101",
				"101010111101",
				"101010111101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"011111011101",
				"011111011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001100",
				"011110111100",
				"011110111011",
				"011010011010",
				"010001110111",
				"001000110011",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000110011",
				"001101110111",
				"011010111011",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100111011111",
				"100111011111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"101011101111",
				"101011011111",
				"101011001110",
				"101011001110",
				"101011001110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100111011110",
				"101011011110",
				"100111001110",
				"100111001101",
				"101011011110",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101011101110",
				"101011101111",
				"100111011110",
				"100111011110",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111111111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111001101",
				"101010111101",
				"101010101100",
				"100110011011",
				"101010101100",
				"101111001110",
				"101111101111",
				"101011101111",
				"100011011101",
				"011111001101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110101011",
				"100010111100",
				"100111011110",
				"100111011101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011111001100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010001001",
				"010101111000",
				"010101100111",
				"011010001001",
				"100010111100",
				"100111001100",
				"011110111100",
				"011010101010",
				"010110101010",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001100111",
				"001101010110",
				"001101000101",
				"001101010110",
				"010101111000",
				"011010001001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010110001000",
				"100111001100",
				"110111101111",
				"111011101111",
				"110111101111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001100",
				"101111001101",
				"101111001100",
				"101010111011",
				"101110111100",
				"101111001100",
				"110011001101",
				"110111011101",
				"111011101110",
				"110111011101",
				"110111011100",
				"110011011100",
				"110011011101",
				"110011011100",
				"110011001100",
				"110011011100",
				"110011011100",
				"110011011100",
				"110011011100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101001",
				"100110001000",
				"101010011001",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"101110111011",
				"101010101011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100110011001",
				"101010111010",
				"110011001100",
				"110011011100",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011101",
				"110111011100",
				"110111011100",
				"110111011100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010111010",
				"101010111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110101001",
				"100010101001",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"101010111011",
				"100110111011",
				"100110101010",
				"100010101010",
				"100010011001",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100010101011",
				"100110111011",
				"100010111011",
				"100110101011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111011",
				"101110111100",
				"101111001100",
				"101110111100",
				"101010111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001100",
				"011110111100",
				"011110101011",
				"010110001001",
				"001101010110",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000101000100",
				"010010001000",
				"011110111100",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111101111",
				"101011011111",
				"100111001110",
				"100110111101",
				"101011001101",
				"101111011110",
				"101111101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011011110",
				"101011011111",
				"101011101111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100011111111",
				"100011101111",
				"100111101111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101011001110",
				"100110111100",
				"100110111100",
				"101111011110",
				"110011111111",
				"101111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100010111100",
				"100111001101",
				"100010111101",
				"100010111101",
				"100010111100",
				"100010101011",
				"100010101011",
				"100110101100",
				"100110011011",
				"100110011011",
				"101111001101",
				"110011101111",
				"101011011110",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110011010",
				"011110001001",
				"100010011010",
				"011110001001",
				"011001111000",
				"011010011010",
				"100011001100",
				"100111011101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110011010",
				"011010001001",
				"011001111000",
				"011001111000",
				"011110011010",
				"100010101011",
				"100010111100",
				"011110111100",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001100110",
				"001101010110",
				"010001100111",
				"010101111000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"101011001100",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110111001101",
				"110111011110",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010101010",
				"101010011001",
				"100110001000",
				"100110001000",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101010111011",
				"101010101010",
				"101110111011",
				"101111001100",
				"101110111011",
				"101010101010",
				"100110101010",
				"100110011001",
				"100110011001",
				"100110101001",
				"101010101010",
				"101110111011",
				"110011001100",
				"110011001100",
				"110111011100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011100",
				"110111011101",
				"110111011100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101001",
				"101010101001",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100010011001",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100010101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100010101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101010111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100011001100",
				"100111001101",
				"100111011101",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111001101",
				"011011001101",
				"011011001100",
				"011110111100",
				"011110101011",
				"010101111000",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001001010101",
				"010110011010",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100111101111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111101111",
				"100111011111",
				"100111001110",
				"100110111101",
				"101011001110",
				"101111011110",
				"101111101111",
				"101111111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011101110",
				"100011101110",
				"100111101110",
				"100011101110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101011001101",
				"101010111101",
				"101110111101",
				"100110011011",
				"100010011010",
				"100110111100",
				"101111011110",
				"101111111111",
				"100111111111",
				"100011101110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"100010101100",
				"011110011011",
				"100010011011",
				"101010101100",
				"101110101100",
				"110011001110",
				"110011011110",
				"101011011110",
				"100111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011101",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"011111001101",
				"100011001101",
				"011111001100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010001001",
				"011110001001",
				"100001111001",
				"011101111000",
				"011010001000",
				"011110101011",
				"100111011110",
				"100111011110",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010001001",
				"011001111000",
				"011001111000",
				"011110001001",
				"100111001100",
				"100010111100",
				"011110111011",
				"011010101010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010101111000",
				"010001100111",
				"010001100111",
				"010101110111",
				"011010001001",
				"011010011010",
				"011010011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110001001",
				"010001110111",
				"011010001001",
				"101011001101",
				"110011101110",
				"111011111111",
				"111011111111",
				"110111101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"111011101110",
				"110111101110",
				"110111101110",
				"110111101110",
				"110011011101",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011001100",
				"101111001100",
				"101110111011",
				"110011011101",
				"110111101110",
				"110111101110",
				"110011011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010101001",
				"101010011001",
				"100110001000",
				"100110001000",
				"101110101010",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111011",
				"101010101010",
				"101010111011",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010111010",
				"101110111010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101110111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111011100",
				"110011001100",
				"110011001011",
				"110011001100",
				"110111011101",
				"110111011100",
				"110011001011",
				"110010111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101010101001",
				"100110011000",
				"100110011000",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101010",
				"101010111010",
				"101110111011",
				"101010111010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111010",
				"101010111010",
				"101110111010",
				"101010111010",
				"101010111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110101010",
				"100110101010",
				"101010101011",
				"101010101010",
				"101010111010",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010101010",
				"100110101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100010101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110101011",
				"100110101011",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111011",
				"101010111011",
				"101010111011",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010101011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100110101011",
				"100110111011",
				"100110111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111011110",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111011",
				"011010011010",
				"010001100111",
				"000100100011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000110011",
				"001101110111",
				"011010101011",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111011111",
				"100111011110",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111101111",
				"100111011110",
				"100111001110",
				"101011001110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100111011110",
				"100111001101",
				"100110111101",
				"101010101100",
				"101010101100",
				"100110001010",
				"101010011011",
				"110011001110",
				"110011101111",
				"101011111111",
				"100011111111",
				"100011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100011001101",
				"100010111100",
				"100010101011",
				"100110011011",
				"101010011100",
				"110010111101",
				"110111011111",
				"110011011111",
				"101011011110",
				"100011011101",
				"011111011101",
				"011111011101",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010001010",
				"100010001001",
				"011101111000",
				"011001111000",
				"011110011010",
				"100111001100",
				"100111011101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011011001100",
				"011010111011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010001001",
				"011010001001",
				"010101111000",
				"010101101000",
				"011001111000",
				"011110001001",
				"100110101011",
				"100010111100",
				"011110111011",
				"011010101011",
				"010110101010",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101111000",
				"010101111000",
				"011010001001",
				"011110011010",
				"011110101010",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"011110011010",
				"100110111011",
				"110011101110",
				"111011111111",
				"111011101111",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111101110",
				"111011101110",
				"111011101110",
				"110111101110",
				"110011011101",
				"110011001100",
				"101111001100",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101111001011",
				"110111011101",
				"110111101101",
				"110111011101",
				"110111011110",
				"111011011110",
				"111011011110",
				"110111011110",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"101110111011",
				"101110101010",
				"101110101001",
				"101010011000",
				"100110001000",
				"101010011001",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111011",
				"101110111010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101110111010",
				"101010101010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101010101001",
				"101010101010",
				"101010011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"110011001100",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110111011100",
				"110011001011",
				"101110111010",
				"101110111010",
				"110011001011",
				"110010111011",
				"101110101010",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101010111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010111011",
				"101110111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110101010",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010101011",
				"101010101010",
				"101010101011",
				"101010111011",
				"101110111011",
				"101010101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"101010111010",
				"101010111011",
				"101010111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101011",
				"101110101011",
				"101110111011",
				"101010111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"101010101011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110101011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"011110011001",
				"011110011001",
				"011110011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100110111100",
				"101010111100",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111011101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011010101011",
				"010110001001",
				"001101010101",
				"000000010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001000100",
				"010110001001",
				"011110111100",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"011111001101",
				"100011011101",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100011111111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011101111",
				"100111101111",
				"100111011111",
				"100111011110",
				"100111011110",
				"101011011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111101111",
				"100111011111",
				"101011011111",
				"101111101111",
				"110011101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101111011111",
				"110111111111",
				"110011111111",
				"101111101111",
				"101011101110",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100111101110",
				"100111011101",
				"101010111101",
				"101010101100",
				"101010011011",
				"110010111101",
				"111011101111",
				"110011111111",
				"101011101111",
				"100111101110",
				"100111111111",
				"100111111111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100010111100",
				"100010101011",
				"100010001010",
				"100110001010",
				"101110101100",
				"110111011111",
				"110011101111",
				"101011101110",
				"100011011101",
				"011111011101",
				"011111101110",
				"100011101110",
				"100011101110",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110011010",
				"100010001001",
				"011101111000",
				"011101111000",
				"100110111011",
				"101011011101",
				"100011001101",
				"011110111100",
				"011111001101",
				"100010111101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011011001100",
				"010111001100",
				"010111001011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010001001",
				"010101111000",
				"010101100111",
				"010101111000",
				"100010001001",
				"100110101011",
				"101010111100",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110001001",
				"010101111000",
				"010101110111",
				"010101111000",
				"011010001001",
				"011110011010",
				"011110011010",
				"011010011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001000",
				"010110001001",
				"010110001001",
				"011010001001",
				"100010101010",
				"110011101110",
				"111011111111",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111101111",
				"111011101110",
				"111011101110",
				"110111011101",
				"110011001100",
				"110010111100",
				"110010111011",
				"110111001100",
				"110111011101",
				"110111001100",
				"110010111011",
				"101110111011",
				"110011001100",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101110111011",
				"101110111010",
				"101010101001",
				"101010101001",
				"100110000111",
				"011101100101",
				"100001110110",
				"101110101010",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010011001",
				"100110011001",
				"101010011001",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"110011001011",
				"110111001100",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001011",
				"101110111010",
				"101110111010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101010111010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010101010",
				"100110101010",
				"100110011001",
				"100010011010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"100110101010",
				"100110011001",
				"100110011001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110011001",
				"100010011001",
				"100110101010",
				"100010101001",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"100110101011",
				"100010101010",
				"100010011010",
				"100010101010",
				"100010011010",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011010111011",
				"010110011010",
				"010001110111",
				"000100110100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001001010110",
				"011010101010",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101110",
				"100111101110",
				"100111101110",
				"101011101110",
				"101011101110",
				"101011011110",
				"100111001101",
				"100110111100",
				"101010111101",
				"101111011110",
				"110011111111",
				"110011111111",
				"101111101111",
				"101011101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011111111",
				"100111101111",
				"100111011110",
				"101011001101",
				"101110111100",
				"101110101100",
				"110010111101",
				"111011101111",
				"110011101111",
				"101111101110",
				"101011101110",
				"100111101110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"011111011110",
				"011111011110",
				"011111011101",
				"100011011110",
				"100011001101",
				"100010111101",
				"100110111101",
				"100110011011",
				"100110001010",
				"110010111101",
				"111011101111",
				"101111011110",
				"100111011101",
				"100011011101",
				"100011101110",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111011101",
				"011111001101",
				"011111011101",
				"011111001101",
				"011110111100",
				"011010111011",
				"011110101011",
				"011110101011",
				"011110011011",
				"011101111001",
				"100001111000",
				"100010011010",
				"101011001101",
				"101011011110",
				"100011001101",
				"011110111100",
				"100011001101",
				"100011001101",
				"100010111101",
				"100010111100",
				"011110111100",
				"011110111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011110011010",
				"011001111001",
				"010101100111",
				"011001111000",
				"100110101011",
				"101010111100",
				"100110111011",
				"011110111011",
				"011010111011",
				"010110101010",
				"010110111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110001001",
				"010010001000",
				"010010001000",
				"010110001000",
				"010101111000",
				"010001100111",
				"001101010110",
				"010001100110",
				"010101111000",
				"011110011010",
				"011110011010",
				"011010011001",
				"010110001001",
				"010110011001",
				"010010001000",
				"001110001000",
				"010110011001",
				"010010001000",
				"001101110111",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001000",
				"010101110111",
				"100110101011",
				"110111101110",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"110111001100",
				"110011001100",
				"110111011101",
				"111011101110",
				"111011011101",
				"110011001100",
				"110011001100",
				"110111011101",
				"110111011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110010111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"110011001011",
				"101110111010",
				"101010101010",
				"101010101001",
				"100001110111",
				"010101000100",
				"011001010100",
				"101010011000",
				"110010111011",
				"101110111011",
				"110010111011",
				"101110111011",
				"101010111010",
				"101010111011",
				"101111001100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101001",
				"101010101010",
				"101010101010",
				"101110111010",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110011001",
				"100110011000",
				"101010011001",
				"101110101010",
				"110010111011",
				"110011001011",
				"110010111011",
				"101110101010",
				"101110101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"100110101001",
				"100010011001",
				"100010011001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"100110011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010101010",
				"100110011001",
				"100010011000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100010011000",
				"100010011000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"101010101011",
				"101010101011",
				"100110101011",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010101010",
				"100110101010",
				"100110111011",
				"100110101011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"100110111101",
				"100111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111011",
				"010110011001",
				"001101010110",
				"000100100011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000110011",
				"010010001000",
				"011010111011",
				"011111001101",
				"100011011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"100111101111",
				"100111101110",
				"100111101110",
				"100111011110",
				"100111001101",
				"100110111101",
				"101010111101",
				"110011001110",
				"110111101111",
				"110011111111",
				"101111111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111001101",
				"101010111101",
				"101010101100",
				"110011001110",
				"111111111111",
				"111011111111",
				"110011101110",
				"101111101110",
				"101011101110",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100111001101",
				"100010101100",
				"100010011011",
				"101010101100",
				"101111001101",
				"110111101111",
				"110011011111",
				"101111011110",
				"100111011110",
				"100111011101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011101",
				"100011011101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011101",
				"100011011101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010101011",
				"100010001010",
				"100001111001",
				"100010011010",
				"101010111100",
				"101111011110",
				"101011001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011110011011",
				"011110001010",
				"011001111000",
				"010101100111",
				"011110001001",
				"100110111100",
				"100110111100",
				"011110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010101111000",
				"010101100111",
				"010001010110",
				"010001010110",
				"010101100111",
				"011010001001",
				"011110101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010110001000",
				"010101110111",
				"011010001000",
				"101111001101",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"111011101110",
				"111011101110",
				"110111101110",
				"110111011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"110011001011",
				"101111001011",
				"101111001011",
				"101110111010",
				"101010011001",
				"100110011000",
				"100110001000",
				"100110000111",
				"011101100110",
				"100001110111",
				"101010101001",
				"101110111011",
				"101110111011",
				"101010101010",
				"101010111011",
				"101010111011",
				"101111001100",
				"101111001100",
				"101011001100",
				"101010111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010101010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110011001",
				"100010001000",
				"100010000111",
				"101010011001",
				"101010101001",
				"101110101010",
				"101110111010",
				"101110101001",
				"101010101001",
				"100110011000",
				"100110011000",
				"100110001000",
				"101010101001",
				"101110111010",
				"101010101001",
				"100110011000",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"100110101001",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110011001",
				"100010011000",
				"100010011000",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011010",
				"101010011001",
				"100110011001",
				"100010001000",
				"100010001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100110011001",
				"100110101001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110001000",
				"011110001000",
				"100010011001",
				"100010011000",
				"100010011001",
				"100010011001",
				"100010011010",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100010101011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"100110111101",
				"100110111101",
				"100111001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111011",
				"011110101010",
				"010110001000",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001010101",
				"010110011001",
				"011010111100",
				"011111001101",
				"100011011110",
				"011111001110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111011110",
				"101011011110",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011011110",
				"101011001110",
				"101111001101",
				"110111011110",
				"111011111111",
				"110011111111",
				"101111111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111001110",
				"100110111101",
				"101010111101",
				"110011001110",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011111111",
				"101111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111001110",
				"100111001101",
				"100010101100",
				"011110011010",
				"100110101011",
				"101111001101",
				"111011101111",
				"110111101111",
				"110011011111",
				"101111011110",
				"101011011110",
				"100111011110",
				"100011011101",
				"100011011101",
				"100011011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010101011",
				"011110001010",
				"011101111001",
				"100010001010",
				"100110101100",
				"101111001110",
				"101111011110",
				"101011001101",
				"100111001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011110101011",
				"011110101011",
				"011110001010",
				"011001101000",
				"011001101000",
				"100010011010",
				"100110111100",
				"100110111100",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110001001",
				"010101111000",
				"010101100111",
				"010101000110",
				"010101010110",
				"011001111000",
				"011110011010",
				"011110101011",
				"011010101010",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010001111000",
				"010101111000",
				"010101110111",
				"010001100110",
				"011010001000",
				"101110111100",
				"110111011110",
				"111111111111",
				"111011101111",
				"111011101110",
				"111011101110",
				"111111111111",
				"111111111111",
				"111111101111",
				"111111101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011101111",
				"110111101110",
				"110011011101",
				"110111011110",
				"110111011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101111001011",
				"101110111011",
				"101110111010",
				"101010111010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101111001011",
				"101111001011",
				"101110111010",
				"101110111010",
				"101010101001",
				"101010011000",
				"101010011000",
				"100110011000",
				"100010000111",
				"100110001000",
				"101010011001",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010101010",
				"100110011001",
				"100010011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"100110011001",
				"100110011000",
				"100010001000",
				"100110011001",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010101001",
				"101010011001",
				"100110011000",
				"100110011000",
				"101010101001",
				"101010101010",
				"100110101001",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100010011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110101001",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011001",
				"100010001000",
				"011110000111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110001000",
				"100010000111",
				"011110000111",
				"100010001000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100010000111",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010001000",
				"100010001000",
				"011101110111",
				"011001110111",
				"011001110111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011000",
				"100010011000",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100110111100",
				"100110111101",
				"100111001101",
				"100111001100",
				"100011001100",
				"011110111011",
				"011110101011",
				"011010011001",
				"010101110111",
				"001000110011",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001101100110",
				"011010101010",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011110",
				"011111011111",
				"011111011111",
				"100011011110",
				"100011011111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111011110",
				"101011101111",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011011110",
				"101111001101",
				"110111011110",
				"111011111111",
				"110111111111",
				"110011111111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111011111",
				"100111001110",
				"100110111100",
				"101111001110",
				"110111101111",
				"111111111111",
				"111011111111",
				"110111101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100111001101",
				"100010101100",
				"011110011010",
				"100110101100",
				"110011011110",
				"110111101111",
				"110111101111",
				"110011011111",
				"101111011111",
				"101111101111",
				"101011011110",
				"100111011110",
				"100111011101",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010101011",
				"100010001010",
				"011101111001",
				"011110001001",
				"101010111100",
				"110011011110",
				"101111011110",
				"101011011110",
				"101011011101",
				"100111001101",
				"100111001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110101011",
				"011110001010",
				"011001111000",
				"011001111000",
				"100010011010",
				"101010111100",
				"100110111100",
				"100010111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010101010",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010101100111",
				"010101010110",
				"011001111000",
				"100010011010",
				"100010101011",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010001111000",
				"010001110111",
				"010001100111",
				"001101010110",
				"010001010110",
				"011101111000",
				"100110011010",
				"101110111011",
				"110011011101",
				"110111101110",
				"110111101110",
				"110111101110",
				"111011101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101111",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011001100",
				"101110111100",
				"101110111011",
				"110011001011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101001",
				"100110101001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110011000",
				"100110011000",
				"101010011001",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110011001",
				"100110101001",
				"100110011001",
				"100010001000",
				"100010000111",
				"100010000111",
				"100110011000",
				"101010101001",
				"101110101010",
				"101110111010",
				"101110101001",
				"101010101001",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010101001",
				"101010011000",
				"100110011000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010000111",
				"100010000111",
				"011110000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100010000111",
				"100010000111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"011110000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"011101110111",
				"011001100110",
				"011001100110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110000111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010000111",
				"011101110110",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110111",
				"011001110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010011000",
				"100010001000",
				"011110001000",
				"011110000111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100010111100",
				"100010111011",
				"011110101010",
				"011010011001",
				"010001100110",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100110",
				"011010101011",
				"011111001101",
				"011111011110",
				"100011011111",
				"100011011110",
				"011111011111",
				"011111011110",
				"011111011111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"110011111111",
				"110011111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111101111",
				"101011011101",
				"101011001100",
				"110011011110",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111101111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111011110",
				"100111001110",
				"100110111100",
				"110011011111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100111011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010101100",
				"101011001101",
				"110111101111",
				"110111101111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111011",
				"011110111011",
				"011110111100",
				"100010101100",
				"100010011010",
				"011101111001",
				"100010011010",
				"101111001101",
				"110011011110",
				"101111001101",
				"101011001101",
				"101011011101",
				"100111011101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100011001100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011110101011",
				"011110011010",
				"011001111001",
				"011001111000",
				"100010001010",
				"101010111100",
				"101011001101",
				"100111001100",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010101100111",
				"011001100111",
				"011110001001",
				"100010101011",
				"100010101011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010001111000",
				"010001111000",
				"010001100111",
				"001101010110",
				"010001100111",
				"011001111000",
				"011001110111",
				"011001111000",
				"100110101010",
				"101111001100",
				"110111011110",
				"110111101110",
				"111011101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111101111",
				"111011101111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101110",
				"110111001101",
				"110111001101",
				"110111011101",
				"110111011101",
				"111011101110",
				"110111011101",
				"110011001100",
				"101110111011",
				"101110111010",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"100110101001",
				"100110101001",
				"101010101001",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010011000",
				"101010101001",
				"101110111011",
				"101110111011",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010011000",
				"100010001000",
				"100010001000",
				"100110011001",
				"101010101001",
				"101010011001",
				"101010011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"100110101001",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010101001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100001110111",
				"011101110110",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100001110111",
				"011101110110",
				"011101110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110110",
				"011001100110",
				"010101100101",
				"010101100101",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001100110",
				"011001110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011001100110",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001100110",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101100110",
				"011001100110",
				"011001110110",
				"011001110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"100010001000",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011010",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110101010",
				"010110001000",
				"001101010101",
				"000000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101100111",
				"011010101011",
				"011111001101",
				"011111011110",
				"100011011110",
				"011111011110",
				"011111011111",
				"011111011110",
				"011111011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111001110",
				"101011001101",
				"101111011110",
				"110111111111",
				"110011101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"100111001101",
				"100111001100",
				"110011011110",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101110",
				"100011101111",
				"100111101111",
				"100111011110",
				"100111001101",
				"100111001101",
				"110011101111",
				"111011111111",
				"110111101111",
				"110011011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011111",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010111100",
				"101011001101",
				"110011011110",
				"110111101111",
				"110011011110",
				"101111001110",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111011101",
				"100111011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001100",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110001001",
				"100010011010",
				"101010101100",
				"110011001101",
				"101111001101",
				"101010111100",
				"100110111100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110101011",
				"011010101010",
				"011010011010",
				"011110001010",
				"011001111001",
				"011001111000",
				"100010001010",
				"101010111100",
				"101111001101",
				"101011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010101100111",
				"011001100111",
				"011101111000",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010001111000",
				"010010001000",
				"010110001000",
				"010001100111",
				"001101010110",
				"010101110111",
				"011110001001",
				"011110001001",
				"011110001000",
				"011010001000",
				"011110011001",
				"101111001100",
				"110111101110",
				"110111101110",
				"110111101110",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111101111",
				"111111111111",
				"111111101111",
				"111011011110",
				"110011001100",
				"101110111011",
				"110111001100",
				"110111001100",
				"110111011101",
				"110111011101",
				"110011001100",
				"101110111011",
				"101110111010",
				"101010101010",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101110111011",
				"101111001100",
				"110011001100",
				"101111001011",
				"101110111011",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101110111010",
				"101010101001",
				"101010011001",
				"101010101001",
				"101010011001",
				"100110011001",
				"101010011001",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011000",
				"100010001000",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100110011001",
				"100110011000",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110101001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"010101100110",
				"010101100110",
				"010101010101",
				"010101100101",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101100110",
				"011101100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"100010011010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011010011001",
				"010001110111",
				"001000110100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"010001110111",
				"011010111011",
				"011111001101",
				"011111011110",
				"100011011110",
				"011111011110",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"110111101111",
				"111011111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"100111011101",
				"101011001101",
				"110011101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111001101",
				"101111011111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001101",
				"100011001101",
				"100011001100",
				"100010111100",
				"100111001101",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001100",
				"101011001101",
				"101111011101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"100111001100",
				"100111001100",
				"100011001100",
				"100010111100",
				"100011001100",
				"100011001100",
				"011110111011",
				"011110101011",
				"011010101011",
				"011110011010",
				"011110001001",
				"101010111100",
				"110011011101",
				"101111001101",
				"101011001100",
				"101011001100",
				"100111001100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100010111100",
				"100010111100",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010001001",
				"011001111000",
				"011101111001",
				"100110101011",
				"101111001101",
				"101011001100",
				"100110101011",
				"100010111011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010101100111",
				"010101100111",
				"011001111000",
				"100010101011",
				"100110111100",
				"100010111011",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001100111",
				"001101010110",
				"010101110111",
				"011110011010",
				"100010101010",
				"011010001001",
				"011010001000",
				"011010001000",
				"011110011001",
				"101010111100",
				"110011101110",
				"110111101111",
				"110111101110",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101110",
				"110111011101",
				"110010111100",
				"110010111100",
				"110010111100",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110011001100",
				"110011001011",
				"101111001011",
				"110011001100",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101111001011",
				"101110111011",
				"101010111011",
				"101010111010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"100110011001",
				"100110011001",
				"101010111010",
				"101010111010",
				"101110111010",
				"101110111010",
				"101010101001",
				"100110011000",
				"100110011001",
				"101010011001",
				"100110011001",
				"101010101010",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101010",
				"101010111010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100010011001",
				"100010001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100001110111",
				"011101110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110110",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010101100101",
				"010101100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011001110110",
				"011001100110",
				"011001100110",
				"010101100101",
				"010101010101",
				"010101010110",
				"010101010110",
				"010101010110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101100110",
				"011101100110",
				"011101100110",
				"011101100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011001110111",
				"011001111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011010001000",
				"001101010101",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111011",
				"011111011101",
				"100011011110",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011101111",
				"110111111111",
				"111011111111",
				"110011101111",
				"110011101110",
				"110011101110",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101011011101",
				"101111101110",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111001110",
				"100111001110",
				"110011101111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101111011111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101111011110",
				"110011101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001100",
				"100011001100",
				"100010111100",
				"100111001100",
				"101011001100",
				"101011001101",
				"101111011101",
				"101111011110",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100010111100",
				"100011001100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110011010",
				"100110101011",
				"101111001101",
				"110011011110",
				"101111001101",
				"101010111100",
				"101011001100",
				"100111001100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100111001100",
				"100111001100",
				"101011001101",
				"100111001100",
				"100110111100",
				"100010111011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011110011010",
				"011110011010",
				"011010001001",
				"011110001001",
				"100010011010",
				"101010111100",
				"101011001101",
				"100110111100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010101110111",
				"011001111000",
				"011110001001",
				"100110101011",
				"100110111100",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110001001",
				"010001111000",
				"010001100111",
				"010001100111",
				"011010001000",
				"011110011010",
				"011110011010",
				"011010001001",
				"011110011001",
				"011010011001",
				"010110001000",
				"011010001001",
				"100110111011",
				"101111011101",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001100",
				"110010111100",
				"110011001100",
				"111011011101",
				"111011011101",
				"110111011101",
				"110111011101",
				"110111011100",
				"110011011100",
				"110011011100",
				"110011011100",
				"110011011100",
				"101010111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101111001100",
				"101111001100",
				"101111001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110101001",
				"101010101010",
				"101111001011",
				"101111001011",
				"101010111010",
				"101010101010",
				"101010101001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101110111011",
				"101110111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100010011001",
				"100010011001",
				"100110101001",
				"100110101010",
				"101010101010",
				"101010111011",
				"100110101010",
				"100110101010",
				"100010101001",
				"100010011001",
				"011110011000",
				"011110001000",
				"011010000111",
				"011001110111",
				"011001110111",
				"011110000111",
				"011110001000",
				"011110000111",
				"011101110111",
				"011110000111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011101110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011101111000",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110110",
				"011001110111",
				"011001110110",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001100111",
				"011001100111",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011101111000",
				"011001111000",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001100111",
				"011001100111",
				"011001110111",
				"011001110111",
				"011001100110",
				"011001100110",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001001",
				"011110001001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"011110011010",
				"100010011010",
				"100010101010",
				"100010101010",
				"011110011001",
				"010101110111",
				"001001000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001001100110",
				"011010101011",
				"011111011110",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"100011101111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011101110",
				"101011111111",
				"101111111111",
				"101111101110",
				"110011111111",
				"111011111111",
				"111011111111",
				"110011101111",
				"110011101110",
				"101111101110",
				"101111101110",
				"101111101111",
				"101111101111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101111011111",
				"110011111111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101111101111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111011110",
				"110011101111",
				"110111101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001100",
				"100011001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"101011001100",
				"101011001101",
				"101011011101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010101011",
				"100010111011",
				"100110111100",
				"100110111100",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001100",
				"100111001100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100010111011",
				"100010111011",
				"011110101011",
				"100010111011",
				"100010111011",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001100",
				"100010111100",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"100010011010",
				"100010011010",
				"011110001001",
				"100010011010",
				"100110111100",
				"101011001100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101010",
				"100010111011",
				"100110111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"011010101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001000",
				"010101111000",
				"011110001001",
				"100110101011",
				"100110111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010111011",
				"011110101011",
				"011110101011",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001100111",
				"010001100111",
				"011010011001",
				"100010101011",
				"011110101010",
				"011110101010",
				"011010011001",
				"011010001001",
				"011010011001",
				"010110001000",
				"011010001000",
				"100010101010",
				"101011001101",
				"101011001100",
				"101011001100",
				"101111001100",
				"110011011101",
				"110111011101",
				"110111011101",
				"110011001101",
				"110111011101",
				"110111011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011011100",
				"101111001100",
				"101111001011",
				"101011001011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"100110111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101111001011",
				"101010111011",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101111001011",
				"101010111010",
				"101110101010",
				"101010101001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110011000",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100010101001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011010001000",
				"011110001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011001110111",
				"011001110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"011001111000",
				"011001110111",
				"011001110111",
				"011001111000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"011001110111",
				"011001110111",
				"011001111000",
				"011001111000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011110001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011110001000",
				"011101111000",
				"011101111000",
				"011101111000",
				"011101111000",
				"011001110111",
				"011001110111",
				"011001110111",
				"011010000111",
				"011010001000",
				"011110011001",
				"100010011010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010011010",
				"011110011001",
				"011110001001",
				"011110001001",
				"011010001000",
				"011001111000",
				"011010001000",
				"011110001000",
				"011110001000",
				"011101110111",
				"011001110111",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001010101",
				"011001010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011101110110",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001001",
				"100010001001",
				"100010001001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"100010011010",
				"011110011010",
				"011010001000",
				"010001100110",
				"001000100011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101100111",
				"010110101011",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100011101111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011101110",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111101110",
				"110011101111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011101111",
				"101111101111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101111011110",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111001101",
				"101111001101",
				"110011011110",
				"110111101111",
				"110111101111",
				"110011101111",
				"101111011110",
				"101111011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"100110111100",
				"101010111100",
				"101011001101",
				"101111001101",
				"101111011110",
				"101011001101",
				"101011001100",
				"100110111100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100011001100",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100111001100",
				"101011001101",
				"101011001101",
				"100110111100",
				"100010101011",
				"100110101011",
				"100110101011",
				"100110011011",
				"100110011010",
				"100110011010",
				"100110101011",
				"101011001100",
				"100111001100",
				"100010111011",
				"011110111011",
				"100011001100",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010111011",
				"100010111100",
				"100010111100",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010101111000",
				"011001111000",
				"100010011010",
				"100110111011",
				"100010101011",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110111011",
				"011110111011",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010001111000",
				"010001110111",
				"010110001000",
				"011110011010",
				"011110101011",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011110011001",
				"101010111011",
				"110011011101",
				"110111011110",
				"110011011101",
				"110011011101",
				"111011101110",
				"110011011101",
				"101111001100",
				"101111001011",
				"101011001011",
				"101011001011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100010011001",
				"100110101001",
				"100110011001",
				"100010011001",
				"100110101001",
				"100110101010",
				"100110101010",
				"101010101010",
				"100110101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100010000111",
				"011101110111",
				"011110000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010001000",
				"100010011000",
				"100110011001",
				"100110011001",
				"100010011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101100111",
				"010101110111",
				"011010001000",
				"011010001001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101110111",
				"010101111000",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010001001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010101011",
				"011110101011",
				"100010101011",
				"100010011010",
				"011110011010",
				"100010011010",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010101010",
				"100110101011",
				"100110111100",
				"101011001101",
				"101011001100",
				"101010111100",
				"101011001101",
				"101011001101",
				"100110111100",
				"100110111100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"100010011001",
				"100010011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011001110111",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001001",
				"011110001001",
				"100010001001",
				"100010011001",
				"011110011001",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110001001",
				"011001110111",
				"001101000101",
				"000100010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100011",
				"001101111000",
				"011010111011",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110111101111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111110",
				"101011101110",
				"101111101110",
				"110011101111",
				"110111111111",
				"111011111111",
				"110111101111",
				"110011101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"110011011111",
				"110111101111",
				"110111111111",
				"110011101111",
				"101111101111",
				"101011011110",
				"101011101110",
				"101011101110",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011011110",
				"101011011110",
				"101111011101",
				"101111011110",
				"110011011110",
				"110011011110",
				"101111001101",
				"101110111100",
				"110011001101",
				"110011011110",
				"110111101111",
				"110111101111",
				"110011011110",
				"101111011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111011101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001100",
				"101010111100",
				"101010111100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101010111100",
				"101110111100",
				"101111001101",
				"101111001101",
				"101111011101",
				"101011001101",
				"100111001100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111100",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010101011",
				"101010101011",
				"100110011010",
				"101010011011",
				"101010101011",
				"101010111100",
				"101011001100",
				"100110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011010001001",
				"011010001001",
				"011010001001",
				"011110001001",
				"100010101010",
				"100110101011",
				"100010101011",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110101011",
				"011110101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010001111000",
				"010101111000",
				"011010001001",
				"011110101010",
				"011110101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"010110001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"011110011001",
				"101010111100",
				"101111011101",
				"101111001101",
				"100110101011",
				"100110101010",
				"100010011001",
				"011110011001",
				"011110011001",
				"011010011000",
				"011010001000",
				"010110000111",
				"010101110111",
				"010101100110",
				"010101100111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110011000",
				"011110011001",
				"011110011001",
				"011010011000",
				"010110000111",
				"010110000111",
				"011010001000",
				"011010001000",
				"011110011000",
				"100010011001",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"101111001011",
				"101110111011",
				"101010111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010001000",
				"100010011000",
				"100110011001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110011001",
				"011110011001",
				"011010001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100111",
				"010101111000",
				"010110001000",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100010111100",
				"100011001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100110101011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100010111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100111001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100110111101",
				"100110111100",
				"100010101100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110011011",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011101110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001001",
				"100010011001",
				"011110011001",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110001000",
				"010101100110",
				"001000110011",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100110011",
				"010010001001",
				"011011001100",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101110",
				"101111011110",
				"110011101111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011101110",
				"101011101110",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"101111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011110",
				"110011011110",
				"110111101111",
				"110111101111",
				"110111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011001101",
				"101011001101",
				"101011001100",
				"101011001101",
				"101010111100",
				"101010111100",
				"101010101011",
				"101110101011",
				"110011001101",
				"110111011110",
				"110111011110",
				"110011011110",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100110111100",
				"100110111100",
				"101010111100",
				"101010101011",
				"100110101010",
				"100110011010",
				"101010101011",
				"101110111100",
				"110011001101",
				"110011011110",
				"101011001101",
				"101011001101",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100110101011",
				"100110101011",
				"101010101011",
				"100110011010",
				"100110001010",
				"100110001001",
				"101010101011",
				"101110111100",
				"101111001100",
				"100110111100",
				"100010111011",
				"100010111011",
				"011111001100",
				"011110111011",
				"011110111011",
				"100010111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"100110111100",
				"100010101011",
				"100010101011",
				"100110101011",
				"100010011010",
				"011110001001",
				"011110001001",
				"011110011010",
				"100110101011",
				"100110101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010001111000",
				"010110001000",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"010110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"001101100110",
				"010001100111",
				"011110011001",
				"100010101010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010011000",
				"011010011000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"011010001000",
				"011110001000",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010101010",
				"100110101010",
				"100110111011",
				"101010111011",
				"101010111011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001011",
				"101110111011",
				"101010111011",
				"100110101001",
				"100110011001",
				"100010001000",
				"100010001000",
				"100010011000",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011001110111",
				"010101111000",
				"010001110111",
				"010001111000",
				"010101111000",
				"010101111000",
				"010001110111",
				"010001100111",
				"010001100111",
				"010101111000",
				"010110001000",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100010111100",
				"100010101100",
				"100010111100",
				"100110111100",
				"100110111101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100110111101",
				"100111001101",
				"100110111101",
				"100110111101",
				"100010111100",
				"100010101100",
				"100010101100",
				"100010101100",
				"100010101100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001001",
				"011110011001",
				"100010011001",
				"011110011001",
				"011110001000",
				"011001100111",
				"001101000101",
				"000100010010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000101000100",
				"010010011001",
				"011111001101",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101110",
				"101111101110",
				"110011101111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011101111",
				"110011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011111111",
				"101111111111",
				"101111111110",
				"101011111110",
				"101011111110",
				"101011101110",
				"101111101110",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"101111111111",
				"101011111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"101111001101",
				"110011001110",
				"110111011111",
				"110111101111",
				"110011011111",
				"101111011110",
				"101011011101",
				"100111011101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101011011101",
				"101011001101",
				"101011001100",
				"101010111100",
				"100110101010",
				"100010011010",
				"100110011010",
				"101110101011",
				"110011001101",
				"110111011110",
				"110011011110",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001100",
				"100111001101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010101011",
				"100110011010",
				"100010001001",
				"100010001001",
				"101010101010",
				"101110111100",
				"110011001101",
				"101111001101",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101010",
				"100010011010",
				"100010001001",
				"100001111001",
				"100110001001",
				"100110011010",
				"101010101011",
				"101110111100",
				"101011001100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100011001100",
				"011110111011",
				"011110111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110011010",
				"100010011010",
				"100010011010",
				"100110101011",
				"100110111100",
				"100110111011",
				"100010101011",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"011010001000",
				"011010001000",
				"010001110111",
				"010001110111",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010001110111",
				"001101100110",
				"001101100110",
				"010001110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110011001",
				"011110001001",
				"100010011001",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101001",
				"011110011001",
				"011110001000",
				"010101110111",
				"010101100110",
				"010101100111",
				"011001110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010101111000",
				"010101111000",
				"010110001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011110101100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101100",
				"100010101100",
				"100010101100",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110011010",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011001110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110001000",
				"011001110111",
				"010001010101",
				"001000100011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001010101",
				"010110011010",
				"011111001101",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111101110",
				"110011101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101111",
				"110011101111",
				"101111111111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101010111100",
				"100110101100",
				"101010101100",
				"110010111101",
				"110111011110",
				"110111011111",
				"110011011110",
				"101111011101",
				"101011001101",
				"101011011101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111001101",
				"101010111100",
				"100110011010",
				"100010011010",
				"100110011010",
				"110010111100",
				"110111001101",
				"110111011110",
				"110011001101",
				"101111001100",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001100",
				"100111001100",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101111001100",
				"101010111011",
				"100110011010",
				"100110001001",
				"100110011010",
				"101110111011",
				"110011001100",
				"101111001100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110101010",
				"100010001001",
				"011101111000",
				"100001111001",
				"101010011010",
				"101110111100",
				"101110111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011110011010",
				"100010101011",
				"100110101011",
				"100010011010",
				"011110001001",
				"100010011001",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101001",
				"010110011001",
				"011010101010",
				"011010011010",
				"011110101010",
				"011110101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010001001",
				"010001111000",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010001110111",
				"010101111000",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"011001110111",
				"011001110111",
				"011001110111",
				"011110001000",
				"100010011001",
				"100010011001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011001",
				"011110001000",
				"011001110111",
				"010101110110",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001100110",
				"010101111000",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010101111000",
				"010110001001",
				"011010001001",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011001",
				"011110001001",
				"011110001000",
				"011001110111",
				"010001010110",
				"001000110011",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101010110",
				"011010101011",
				"011111011101",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101011111111",
				"101011101111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011001101",
				"100110111100",
				"100110101011",
				"101010101100",
				"110010111101",
				"110111011110",
				"110111011110",
				"110011001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011101",
				"101111011110",
				"101111011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011011101",
				"101011001101",
				"101111011101",
				"101111001101",
				"101010111100",
				"100110101010",
				"100110101010",
				"101010101011",
				"110011001101",
				"110111011101",
				"110111011101",
				"101111001101",
				"101111001100",
				"101011001100",
				"101011001101",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010101011",
				"101010011010",
				"101010011010",
				"101110101011",
				"110011001100",
				"110011011101",
				"101111001100",
				"101010111011",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110101010",
				"100010001001",
				"011101111000",
				"100110001001",
				"101010101011",
				"101111001100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"100110101011",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110011010",
				"100010011010",
				"011110001001",
				"011001111000",
				"011001111000",
				"100010011001",
				"100110101011",
				"100110111011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110011001",
				"011110101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010011010",
				"011010011001",
				"010110011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010101111000",
				"010001111000",
				"010110001001",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001001",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001010101",
				"010001100110",
				"010101110111",
				"011001110111",
				"011110001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"001101100110",
				"001101010110",
				"010001100111",
				"010101111000",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101111000",
				"010001100111",
				"010001100111",
				"010001100111",
				"010101111000",
				"011010001001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010110001000",
				"011010001001",
				"011010011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"100010111100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111100",
				"100010101100",
				"100010101100",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"010101100110",
				"001101000100",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111100",
				"100011011110",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011101111",
				"101011101110",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101010111100",
				"101110111101",
				"110111001110",
				"110111001110",
				"110111001110",
				"110011001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"101111011101",
				"101111001101",
				"110011001110",
				"110011001110",
				"110011001110",
				"110011001110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001100",
				"101010111011",
				"100110101011",
				"101010101011",
				"101110111011",
				"110111011101",
				"110111011101",
				"110011011101",
				"101111001101",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010101010",
				"101010011010",
				"101010101010",
				"101110111011",
				"110011001100",
				"110011001100",
				"101111001011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110011010",
				"100010001001",
				"100010001001",
				"100110011010",
				"101010111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"100010111011",
				"100110111011",
				"100110111100",
				"101010111100",
				"101010101100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010011010",
				"011110001001",
				"011101111000",
				"011110001001",
				"100110101010",
				"100110111011",
				"100110111011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110101010",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011010",
				"011110011010",
				"011110101010",
				"011010001001",
				"010110001001",
				"010110001001",
				"011010011010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010001010",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010001001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010001001",
				"011010001000",
				"010101110111",
				"010101100110",
				"010101100110",
				"011001110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010001110111",
				"001101100110",
				"001101100111",
				"010001111000",
				"011010001001",
				"011110011010",
				"011110011010",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"010101111000",
				"010001100111",
				"010001100110",
				"010001100110",
				"010101111000",
				"011010001001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110101010",
				"011010011010",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010001110111",
				"010001110111",
				"010110001001",
				"011010011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011010",
				"011110011010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110011011",
				"011110101010",
				"100010101011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"100010111011",
				"100010111100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"100110111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"100010101011",
				"100010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011110001000",
				"011110001000",
				"011001110111",
				"010101110111",
				"010001010101",
				"000100100011",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101110111",
				"011010111100",
				"100011101110",
				"100111111111",
				"100111111111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101110",
				"110011011110",
				"110011011110",
				"110111101111",
				"111011111111",
				"110111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101010111100",
				"101010111100",
				"101110111101",
				"110111001110",
				"110111001110",
				"110111001101",
				"110011001101",
				"101111001101",
				"101111001100",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011001110",
				"110011001110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101010111011",
				"101010111011",
				"101110111011",
				"101111001100",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011001101",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001100",
				"101011001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001100",
				"110011001100",
				"110011001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101110111011",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001011",
				"101011001011",
				"101010111011",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100010011010",
				"100010001001",
				"100110011001",
				"101110111011",
				"101111001100",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111011",
				"101010101100",
				"101010101100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100110111011",
				"100010011010",
				"011110001001",
				"100010001001",
				"100110101011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111010",
				"011110111011",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010001000",
				"011010001001",
				"011110101010",
				"100010101011",
				"100010101010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011010011001",
				"010110011001",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"010101110111",
				"010101100111",
				"010101110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001100111",
				"010001100111",
				"010101111000",
				"011010001001",
				"011010001010",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011001111000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010001001",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101111000",
				"011010001001",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010001000",
				"010101111000",
				"010101111000",
				"010110001000",
				"011010001001",
				"011110011010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"011110011010",
				"011110011010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010101011",
				"100010101011",
				"100110111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100110111011",
				"100110111100",
				"101011001101",
				"101011001101",
				"100110111100",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010011010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011110001000",
				"011101110111",
				"011001110111",
				"010101100110",
				"001101000100",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101110111",
				"011011001100",
				"100011101111",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011111111",
				"110011111111",
				"101111101111",
				"110011101111",
				"101111101110",
				"101111001101",
				"101010111100",
				"101111001101",
				"110111011111",
				"111011101111",
				"110111101111",
				"110011101110",
				"101111101110",
				"101111101110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101010111100",
				"101010111100",
				"101111001101",
				"110011001101",
				"110111011101",
				"110111011101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101110111100",
				"101010111011",
				"101010111011",
				"101110111100",
				"110011001100",
				"110111011101",
				"110111001101",
				"110111001101",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010101010",
				"101110101011",
				"101110111011",
				"110010111011",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"101010101011",
				"100110011010",
				"100010001001",
				"100110011001",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100010101010",
				"011110011001",
				"011110011001",
				"100110101011",
				"101010111100",
				"101010111100",
				"100110101011",
				"100110101011",
				"100110111011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"100010101011",
				"100010011010",
				"011110001001",
				"011001111000",
				"011001110111",
				"011110011001",
				"100010101010",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110011001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011110011010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011010",
				"100010101010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010011001",
				"011110011001",
				"011010011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010001000",
				"011001111000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001001",
				"011001111000",
				"010101110111",
				"010101110111",
				"011001111000",
				"011010001001",
				"011110011001",
				"011110011010",
				"011010001001",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011001111000",
				"010101111000",
				"011010001000",
				"011110011001",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010001001",
				"011010011001",
				"011010011010",
				"011010001001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010011001",
				"011110011010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011110011010",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010011010",
				"100010101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010111011",
				"100110111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101100",
				"100010111100",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100010001001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001100110",
				"010101010101",
				"001101000100",
				"000100100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101110111",
				"011011001100",
				"100011101110",
				"100111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"101111011110",
				"101110111101",
				"110011001110",
				"110111011111",
				"111011101111",
				"110111101111",
				"110011101110",
				"101111101110",
				"101111101110",
				"101111011110",
				"110011011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101111011110",
				"101111001101",
				"101010111100",
				"101010111100",
				"101111001101",
				"110011001101",
				"110111011101",
				"110111011110",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111011101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101110111100",
				"101010111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110111001101",
				"110111001101",
				"110111001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"101010101010",
				"100110011010",
				"100110011001",
				"101010011010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100010101010",
				"100010011010",
				"100010101010",
				"100110111011",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101010",
				"011110011001",
				"011110001000",
				"011110001000",
				"011110001001",
				"100010011010",
				"100110101010",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010001000",
				"011110001001",
				"100010011010",
				"100010101010",
				"100010101010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010001001",
				"011110001001",
				"011110011001",
				"100010101010",
				"100010011010",
				"011110011010",
				"011110011001",
				"011110011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010001001",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010001001",
				"011110001001",
				"011110011001",
				"011010001001",
				"011010011001",
				"011010011010",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011001111000",
				"011001111000",
				"011110001001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"011010001001",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"100010101010",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"100010011010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010111100",
				"100110111100",
				"100010111100",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010111011",
				"100110111100",
				"100010111100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010111011",
				"100110111100",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101100",
				"100110101100",
				"100110101100",
				"100010101011",
				"100010101011",
				"100010011011",
				"100010011010",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"010101010101",
				"010001000100",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101110111",
				"011011001100",
				"100011101110",
				"100111111111",
				"101011111111",
				"101111111111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"101111001110",
				"110111011110",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110011101110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101111001110",
				"101111001101",
				"101010111100",
				"101110111100",
				"101111001101",
				"110011001101",
				"110111011101",
				"110111011110",
				"110111011101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001101",
				"110111001101",
				"110111001101",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110101011",
				"101010101011",
				"100110011010",
				"100110011010",
				"100110011010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101010",
				"100010011010",
				"100110101010",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010011010",
				"011110011001",
				"011110001001",
				"100010011001",
				"100110101010",
				"100110101010",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010001001",
				"011001111000",
				"100010011001",
				"100010011010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010001001",
				"011110001001",
				"011110011001",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010101111000",
				"011001111000",
				"011010001001",
				"011110001001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010001001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010001001",
				"011110001001",
				"011110001001",
				"011110001001",
				"011110001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011110011001",
				"100010011010",
				"100010101010",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010101010",
				"100010101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101011",
				"100010111011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100110111011",
				"100110111100",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011001100110",
				"010101010101",
				"010001000100",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011011001100",
				"100011101111",
				"100111111111",
				"101011111111",
				"101111111111",
				"101111101111",
				"101111111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110011101111",
				"110011011110",
				"110111011111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101110",
				"110011011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001110",
				"101011001110",
				"101111001101",
				"101111001101",
				"101110111100",
				"101110111100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110111011101",
				"110111001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"110010111100",
				"110011001100",
				"110111001101",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110101011",
				"101010101011",
				"100110011010",
				"101010011010",
				"101010101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101011",
				"101010111011",
				"101110111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010011001",
				"100010011001",
				"100110011010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011001",
				"011010001000",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001000",
				"011001111000",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101110111",
				"010101111000",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010011001",
				"010110001000",
				"010110001001",
				"011010001000",
				"011010001001",
				"011010001001",
				"011110001001",
				"011110001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010101010",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110101010",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"100010101011",
				"100110111011",
				"100110111100",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010101011",
				"100010101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100110011010",
				"100010011010",
				"100110011010",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"010101010101",
				"010001000100",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011011001100",
				"100011111111",
				"101011111111",
				"101011111111",
				"101111111111",
				"101111101111",
				"101111111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"110111101110",
				"110011101110",
				"110111101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111101111",
				"110011101111",
				"110011011110",
				"110111011110",
				"111011011111",
				"111011101111",
				"110111101111",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011011110",
				"110011001110",
				"110011001110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101110111100",
				"101110111100",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"101111001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"100110101011",
				"100110101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010011010",
				"100110101010",
				"100110101010",
				"101010101011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010111011",
				"011110101011",
				"011110101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011001",
				"100010011010",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011110001001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001000",
				"010101111000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101111000",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011110011001",
				"011110011010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011110011001",
				"100010011010",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011110011010",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101011",
				"100110101011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100010101011",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011010",
				"100110011001",
				"100110011001",
				"100110011010",
				"100110011010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"010101010101",
				"010001000100",
				"001100110011",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011011001100",
				"100111111111",
				"101011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011101110",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101110",
				"110011101110",
				"110111101110",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110111011110",
				"110111011110",
				"111011011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"110011001100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110101011",
				"100010101010",
				"100010011010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011110001001",
				"011110001001",
				"011110001001",
				"011110011010",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110011001",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101111000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011010",
				"100010011010",
				"011110101010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011110011001",
				"011110011010",
				"100010101010",
				"100010101010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011110011001",
				"011110011010",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"100010101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101010",
				"100010101010",
				"100010011010",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101010100",
				"001100110011",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111100",
				"100111101111",
				"101011111111",
				"101111111111",
				"101111101111",
				"110011111111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110011111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111100",
				"110010111011",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"101010111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101110111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100010101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"100110101011",
				"101010111011",
				"100110111011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110001001",
				"100010011010",
				"100010011010",
				"100010101010",
				"100010011010",
				"011110011010",
				"011110011001",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001000",
				"011010001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010101111000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"011001111000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011110011001",
				"011110011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011010",
				"100010101010",
				"100010101011",
				"100010101010",
				"100010101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010101010",
				"100010101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010011010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010001000100",
				"001000110010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111100",
				"100111101111",
				"101011111111",
				"101111111111",
				"101111101111",
				"110011101111",
				"110011111111",
				"101111111111",
				"101111111111",
				"101111111111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111100",
				"110010111011",
				"110010111100",
				"110011001100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111011",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"101010101010",
				"101010111010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100110101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110001001",
				"011010001000",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010011001",
				"011010001001",
				"011010001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"100010101010",
				"100010101011",
				"100010101010",
				"100010101010",
				"011110011010",
				"100010011010",
				"100010101010",
				"100010011010",
				"011110011010",
				"100010101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110000111",
				"100110000111",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010101010100",
				"001100110011",
				"001000100001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001001010110",
				"011010111011",
				"100011101110",
				"101011111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111111111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111001101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110011001100",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111011",
				"110011001100",
				"110010111100",
				"110010111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010101010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101011",
				"100110101011",
				"101010101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010011010",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110001001",
				"011110001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110001001",
				"011110001001",
				"011110001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010001001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010101010",
				"100010101011",
				"100010101010",
				"011110011010",
				"011110011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110000111",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010101010100",
				"010001000100",
				"001100110011",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001001010110",
				"010110101011",
				"100011011110",
				"101011111111",
				"101011101111",
				"110011101111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110111001101",
				"110111001101",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111100",
				"110011001100",
				"110011001100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"101010101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110001001",
				"011110001001",
				"011110001000",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"100010011001",
				"011110011001",
				"011110001001",
				"011110001001",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001001",
				"011110011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110011010",
				"011110011001",
				"011110011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011001",
				"100010011010",
				"100010101010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110000111",
				"100110000111",
				"100110000111",
				"100110000111",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010001000100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001001010110",
				"011010101011",
				"100011011110",
				"101011111111",
				"101011101111",
				"110011101111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111101111",
				"110111011111",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110111001100",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010111010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010011010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"011110001001",
				"011110001000",
				"011110001001",
				"011110001000",
				"011110001000",
				"011110001001",
				"011110001001",
				"011110001001",
				"011010001000",
				"011110001000",
				"011110001000",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010001001",
				"011110001001",
				"011110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011010001001",
				"011010001001",
				"011110001001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"011110001001",
				"011110011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"100010011001",
				"100010101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100110000111",
				"100110000111",
				"100110000111",
				"100110000111",
				"100110000111",
				"100110001000",
				"100110000111",
				"100110000111",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010001000100",
				"010001000011",
				"001100110010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111011",
				"100011101110",
				"101011111111",
				"101111101111",
				"110011101111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110111010",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101011001100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010111010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100110101001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110001001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110001000",
				"011110001000",
				"011010001000",
				"011110001001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001001",
				"011110001001",
				"011110001000",
				"011110011001",
				"011110001001",
				"011110001000",
				"011110001000",
				"011110001001",
				"100010011001",
				"100010011001",
				"100110011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110101010",
				"100110101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011010",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100110000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010101010101",
				"010001000100",
				"001101000011",
				"001000100010",
				"001000100001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111100",
				"100011101111",
				"101011111111",
				"101111101111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011011110",
				"111011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111011",
				"110010111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111010",
				"110010111010",
				"110010111010",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100010101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010001001",
				"011110011000",
				"011110011001",
				"011110011000",
				"011110011000",
				"011110001000",
				"011110001001",
				"011110001001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010011000",
				"100010011001",
				"100010011001",
				"100010001001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010011001",
				"100010011001",
				"100110011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010001001",
				"011110001000",
				"100010001000",
				"100010011001",
				"100110011001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001110110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010001010100",
				"010001000100",
				"001100110011",
				"001100110010",
				"001000100010",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011111001100",
				"100011101111",
				"101011111111",
				"101111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011011110",
				"111011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"110010111011",
				"110010111010",
				"110010111010",
				"110010111010",
				"110010111010",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010011001",
				"100010011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010011000",
				"100010011000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010011000",
				"100010011001",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001001",
				"100010011001",
				"100010001001",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"100010011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001001",
				"100010001000",
				"100010001001",
				"100110001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101010101",
				"010001010100",
				"010001000100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101110111",
				"011111001100",
				"100111101111",
				"101011111111",
				"101111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110111011111",
				"110111011111",
				"110111011110",
				"110111011110",
				"110111011110",
				"111011011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101010",
				"100110101001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011101111000",
				"011101110111",
				"011101111000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011101111000",
				"011101111000",
				"011110001000",
				"011001110111",
				"011001110111",
				"011010000111",
				"011010001000",
				"011110001000",
				"011110001000",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011101111000",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001001",
				"100110011001",
				"100110001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010011001",
				"100010001000",
				"011110001000",
				"100010001000",
				"100010011000",
				"100010011000",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011001",
				"100010011000",
				"100110011000",
				"100010011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"010101010101",
				"010101010101",
				"010001000100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"010001111000",
				"011111001101",
				"100111101111",
				"101011111111",
				"101111101111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"110010111010",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101111001100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011101110111",
				"011101111000",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011110000111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011110001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010011000",
				"100010011000",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101010101",
				"010101010101",
				"010001000100",
				"010001000011",
				"001000110010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010010",
				"010001111000",
				"011010111100",
				"100111101111",
				"101011111111",
				"101111111111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111111111111",
				"111111111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111001101",
				"110111001100",
				"110111001101",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101010101001",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101001",
				"101110101010",
				"101110111010",
				"110010111010",
				"110010111010",
				"101110111010",
				"110010111010",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"110010111011",
				"110010111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"100110101010",
				"100110101010",
				"101010111010",
				"101010111011",
				"101011001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010011000",
				"100010001000",
				"100010001000",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110001000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100001110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010001000100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010010",
				"001101110111",
				"011010111100",
				"100111101111",
				"101011111111",
				"101111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111111111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110111011101",
				"110111011101",
				"110111001101",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110101001",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101010",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"110010111010",
				"110010111010",
				"110010111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110111010",
				"101010111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010101001",
				"100010101001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011000",
				"011110011000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"100010011000",
				"100010011000",
				"100010011000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011110000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110000111",
				"100010000111",
				"100010000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001110111",
				"011001110111",
				"011001100110",
				"011001100110",
				"011001100111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001010101",
				"010101010101",
				"010101010100",
				"010001000100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100001",
				"000100010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011010111100",
				"100111101111",
				"101011111111",
				"101111101111",
				"110011111111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101001",
				"101110101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101111001011",
				"110011001011",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101010",
				"101010111010",
				"101010111011",
				"101011001011",
				"101011001100",
				"101011001011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011000",
				"100010011000",
				"100010011000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001100110",
				"011101110110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101100110",
				"011101100110",
				"011001100110",
				"011001100101",
				"011001010101",
				"010101010100",
				"010101000100",
				"010001000100",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001001010110",
				"011010101011",
				"100011101110",
				"101011101111",
				"101111101111",
				"110011111111",
				"110111111111",
				"110011111111",
				"110011111111",
				"110011111111",
				"110111101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"100110101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"101111001011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101011001100",
				"101011001100",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011110000111",
				"011110000111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110110",
				"011001110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100101",
				"010101100101",
				"010101100101",
				"011001100110",
				"011001110110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101100110",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101100110",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100001110111",
				"100001110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101100110",
				"011101100110",
				"011001100101",
				"011001010101",
				"010101010101",
				"010101010100",
				"010001000100",
				"010001000011",
				"001100110010",
				"001000100010",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001001000101",
				"011010101011",
				"100111011110",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110011001",
				"100010011001",
				"100110101001",
				"100110011001",
				"100110101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101001",
				"101110111010",
				"101110111010",
				"101110101001",
				"101110101010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101111001100",
				"110011001100",
				"101111001011",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101001",
				"100010101001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101100101",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001010101",
				"011001010101",
				"011001010101",
				"011001010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101000100",
				"010001000100",
				"001100110011",
				"001000100010",
				"001000010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100110100",
				"010110011010",
				"100011011110",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011011110",
				"111011011110",
				"111011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011000",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100010011001",
				"100110011001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011001110111",
				"010101110110",
				"010101110110",
				"011001110111",
				"011110001000",
				"100010101001",
				"101010111010",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110101010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"101010101001",
				"101010101010",
				"101010101001",
				"101010101010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101011001100",
				"101011001011",
				"101011001100",
				"101011001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111011",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010001010100",
				"010001010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110111",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"010001000011",
				"010000110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100100010",
				"001000100001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000100011",
				"010010001000",
				"100011001101",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111001101",
				"110111001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"101010011000",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"100110101010",
				"100010011001",
				"100010011001",
				"011110011000",
				"011110001000",
				"011001110111",
				"011001110111",
				"011110001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"011101111000",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001010101",
				"001101010101",
				"001101010100",
				"001101010101",
				"010001010101",
				"010101110111",
				"011110001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011000",
				"011110011000",
				"011110001000",
				"011110000111",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001100110",
				"100010011000",
				"100110101001",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101011001011",
				"101011001011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010101010101",
				"010101100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101100110",
				"011101100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001100110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001101100111",
				"011110111100",
				"101011101111",
				"101111111111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100010011001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011001110111",
				"010101110111",
				"010001100110",
				"001101010101",
				"010001100110",
				"010101100111",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101010101",
				"010001010101",
				"011001110111",
				"011110001000",
				"100010011001",
				"100010011000",
				"100010011000",
				"100010011000",
				"100110101001",
				"100110101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110001000",
				"011110001000",
				"100010001000",
				"100110011001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010111010",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101110111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111011",
				"101110111011",
				"101111001011",
				"101111001100",
				"101111001100",
				"101111001011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110111010",
				"101010111010",
				"100110111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"011110000111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001010100",
				"010101010100",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101100110",
				"011101100110",
				"011101100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100100010",
				"001000100010",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001001010110",
				"011010101011",
				"100111011110",
				"101111101111",
				"110011101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110111001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"101010011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100010101010",
				"100010011001",
				"011110011001",
				"011110001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"011001110111",
				"011110001000",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"100110101010",
				"100110101001",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010111010",
				"101010111010",
				"100110111010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101001",
				"100010101001",
				"100010101001",
				"100010101001",
				"100010101001",
				"100010101001",
				"100010011001",
				"100010101001",
				"100010101001",
				"100010101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011110000111",
				"011001110111",
				"011101110111",
				"011101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010001010100",
				"010001000100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010101",
				"010101100101",
				"011001100101",
				"011001100101",
				"011001010101",
				"011001010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010001000100",
				"010001000011",
				"001100110011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001001000101",
				"011010011010",
				"100111011110",
				"101011101111",
				"110011101111",
				"110011111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101110",
				"110111101110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110111001101",
				"110011001101",
				"110011001101",
				"110111001101",
				"110111001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100010011001",
				"011110011001",
				"011110001000",
				"011110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001100111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001000100",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010101110110",
				"011010000111",
				"011110001000",
				"011110001000",
				"011110000111",
				"011010000111",
				"011010000111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011010000111",
				"011110001000",
				"100010011001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101001",
				"100010011001",
				"100010101010",
				"100110101010",
				"100110101010",
				"100110111010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100010011001",
				"100010011001",
				"011110011000",
				"011110011000",
				"100010011000",
				"100010101001",
				"100010101001",
				"100010101010",
				"100010011010",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"100010011001",
				"100010011001",
				"100010101001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"100010011001",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011010001000",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101100111",
				"010101100110",
				"010101100110",
				"010101100111",
				"010101100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100110",
				"010101100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010001010100",
				"010101010100",
				"010101010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101100110",
				"011101100110",
				"011001100110",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100110100",
				"010110001001",
				"100111011101",
				"101011101111",
				"101111101111",
				"110011101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"101010011000",
				"101010011000",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010111010",
				"101010111010",
				"101010101011",
				"100110101011",
				"100110101010",
				"100010101010",
				"011110011001",
				"011110001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001001010110",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100110",
				"011001110111",
				"011110001000",
				"011110011000",
				"011110011001",
				"011110011000",
				"011110001000",
				"011110001000",
				"011110001000",
				"011110000111",
				"011010000111",
				"011010000111",
				"011010000111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011110001000",
				"011110011001",
				"100010011001",
				"100010101001",
				"100010011001",
				"100010011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"011110000111",
				"011110000111",
				"011110000111",
				"011001110111",
				"011001110110",
				"010101110110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010101110110",
				"010101110110",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010101",
				"010001010101",
				"010101100110",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"001101000100",
				"001101000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"010001000011",
				"001101000011",
				"001101000011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000011",
				"010000110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010101000100",
				"010101000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"010001000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010101",
				"010101010101",
				"011001010101",
				"011001010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101000100",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010100",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001010101",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101000100",
				"010001000100",
				"010001000011",
				"010001000011",
				"010001000011",
				"010000110011",
				"010000110011",
				"010001000011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001100110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100011",
				"010001111000",
				"100011001101",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011111111",
				"111011111111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100010101010",
				"100010011010",
				"011110011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001001010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010110",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101010110",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001100110",
				"010101110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"010101100101",
				"010101100101",
				"010001010101",
				"010001010100",
				"001101010100",
				"001101000100",
				"001101000100",
				"001001000011",
				"001001000011",
				"001001000011",
				"001001000011",
				"001001000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"000100100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000000010001",
				"000000010001",
				"000100010001",
				"000100100010",
				"001000110011",
				"001100110011",
				"001101000100",
				"001101000100",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"001000110010",
				"001000110010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100010001",
				"000100010001",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100100001",
				"000100100001",
				"000100100010",
				"000100100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110011",
				"001100100011",
				"001100100011",
				"001100100011",
				"001100110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000100",
				"010101000100",
				"010101000100",
				"010101000100",
				"010101000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"010000110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100100010",
				"001000100010",
				"001000100001",
				"001000100001",
				"001000100001",
				"001000100001",
				"001000100001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101100111",
				"011110111100",
				"101011101110",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"111011011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110101010",
				"100010101010",
				"011110011010",
				"011110011001",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010011000",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001001010110",
				"001001010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010110",
				"001101010110",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010100",
				"001001000100",
				"001001000100",
				"001001010100",
				"001101010100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"000100110011",
				"000100110011",
				"000100110010",
				"000100110010",
				"000100110010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000000010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000010000",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"001000010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100100010",
				"001100110010",
				"001100100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110010",
				"001100110011",
				"010000110011",
				"010000110011",
				"010000110011",
				"001100110011",
				"010000110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"010000110011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"001000010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"001001010110",
				"011110111011",
				"100111101110",
				"101011101111",
				"101111101111",
				"110011101111",
				"110111101111",
				"110111111111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010011000",
				"011010011000",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001000101",
				"001001000101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"000100010000",
				"000100010000",
				"000100010000",
				"000100010000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000010001",
				"001000100010",
				"001000010001",
				"001000010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000101000101",
				"011010101011",
				"100111011110",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110011001",
				"100010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"011010001000",
				"011010001000",
				"010110011000",
				"011010011000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001001010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001000101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101010110",
				"001001010110",
				"001001010110",
				"001001010110",
				"001001100110",
				"001001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101100101",
				"001101100101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001000100",
				"001001000101",
				"001001000101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001000110011",
				"001100110010",
				"001000110010",
				"001000110010",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000101000100",
				"011010101010",
				"100111011110",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"100110011000",
				"101010011000",
				"101010011000",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110011010",
				"100010011001",
				"100010011010",
				"100010011010",
				"011110011010",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001001010110",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000101",
				"001101000101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000110010",
				"001000110011",
				"001000110011",
				"001000100011",
				"000100100010",
				"000100010010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100110011",
				"011010001001",
				"101011011101",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011011111",
				"110111101111",
				"110111101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"101010011000",
				"101010011000",
				"101010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011000",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011001",
				"100010011001",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001101000011",
				"001101000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100011",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"010101110111",
				"100110111100",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111011111",
				"110111101111",
				"111011101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"100110011000",
				"101010011000",
				"101010011000",
				"101010011001",
				"101010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011001",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101100101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001100110100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001101010110",
				"100010101011",
				"101111011110",
				"101111101111",
				"101111101111",
				"110011011111",
				"110111101111",
				"110111101111",
				"111011101111",
				"111011101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"101010011000",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011001",
				"100010011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101010100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001001000100",
				"011110011001",
				"101011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110111011111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011010",
				"100010011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100011",
				"010101110111",
				"100110111100",
				"101111011111",
				"101111101111",
				"110011101111",
				"110011011110",
				"110111011111",
				"110111011111",
				"110111011111",
				"110111011111",
				"110111011111",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001001010110",
				"001001010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101100110",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001101010101",
				"100010101010",
				"101011011110",
				"101111011111",
				"110011101111",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"101010011001",
				"101010011001",
				"101010101001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101010100",
				"001101010100",
				"001101010100",
				"001101010100",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010000",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100110011",
				"011010001000",
				"100110111100",
				"101111011110",
				"110011101111",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100011",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010010",
				"010001100111",
				"100010101011",
				"101111011110",
				"110011101111",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110111001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100101",
				"001101100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110100",
				"011110001001",
				"101111001101",
				"101111011110",
				"110011011110",
				"110111011111",
				"110111011110",
				"110011011110",
				"110011001110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100110",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001000110011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100011",
				"001000100010",
				"000100100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000100010000",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"010101100111",
				"100110111100",
				"101111001101",
				"110011011110",
				"110111101111",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001000100",
				"001101000100",
				"001101000100",
				"001100110100",
				"001100110011",
				"001000110011",
				"001000110011",
				"001100110100",
				"001100110100",
				"001100110100",
				"001100110100",
				"001100110100",
				"001100110011",
				"001000110011",
				"001000110011",
				"001100110011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100100001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000100010000",
				"000100010001",
				"001000010001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"001000100001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000100010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001101000101",
				"011110011010",
				"101011001100",
				"110011011110",
				"110111101111",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011010",
				"100110101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110100",
				"001000110100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001100110011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000100100010",
				"001000100010",
				"001000100010",
				"001000110010",
				"001000110011",
				"001100110011",
				"001000110011",
				"001100110011",
				"001000110010",
				"001000110010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100001",
				"000100010001",
				"001000100001",
				"001000100010",
				"001000110010",
				"001100110010",
				"001100110011",
				"001100110010",
				"001100110010",
				"001000100010",
				"001000100010",
				"001100110010",
				"001100110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000100",
				"001101000011",
				"001100110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100011",
				"010101110111",
				"100110101011",
				"101111001101",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011010",
				"100110011010",
				"100110011010",
				"100110101010",
				"100110011010",
				"100010101010",
				"100010101001",
				"100010011001",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001000110100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"000100100010",
				"000100100010",
				"000100100010",
				"001000100010",
				"001000110010",
				"001000110010",
				"001000110010",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000110010",
				"001000100010",
				"000100100001",
				"001000100001",
				"001000100010",
				"001000100010",
				"001000110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001000100001",
				"000100010001",
				"000100100001",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100110010",
				"001100110011",
				"001100110011",
				"001101000011",
				"001101000011",
				"001101000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100100010",
				"001100100010",
				"001100100010",
				"001000100010",
				"001000010001",
				"000100010001",
				"000100010000",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001101010101",
				"011110011001",
				"101010111100",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110111011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101111000",
				"001101111000",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010101",
				"010001010110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010110",
				"010001010110",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000110010",
				"001000110011",
				"001000110011",
				"001000110011",
				"001100110011",
				"001101000011",
				"001100110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000110010",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"001000100001",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001101000011",
				"010001000100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"001100110011",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100100010",
				"001100100010",
				"001000100010",
				"001000100001",
				"001000100001",
				"001000100001",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000110100",
				"011001111000",
				"100110101010",
				"101111001101",
				"110011011101",
				"110111011110",
				"110111011110",
				"110111011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010110",
				"010001010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000101",
				"001101000101",
				"001101000101",
				"001101000101",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001000110100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110010",
				"000100100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000110010",
				"001100110010",
				"001100110011",
				"001100110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110010",
				"001100110011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001101000011",
				"001100110011",
				"001100110011",
				"001101000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"001101000011",
				"001100110011",
				"010001000011",
				"010001000011",
				"010101000100",
				"010001000011",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100100010",
				"001100110010",
				"001100110010",
				"001000100010",
				"001000110010",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"001000100001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000100010",
				"001101010101",
				"011110001001",
				"101010111011",
				"101111001101",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100110011010",
				"100110011001",
				"100110011001",
				"100110011001",
				"100010011001",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100111",
				"001101100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010110",
				"010001010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001001000011",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000110010",
				"001000110010",
				"001100110011",
				"001101000011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100110011",
				"001101000011",
				"010001000011",
				"010001000100",
				"010001000011",
				"010001000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010101010100",
				"010001000011",
				"010001000011",
				"010001000011",
				"010000110011",
				"001100110010",
				"001100100010",
				"001100110010",
				"001000100001",
				"001000100010",
				"001000110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100110011",
				"010101110111",
				"100010011010",
				"101010111100",
				"101111001101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101110101001",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110011001",
				"100110011001",
				"100110011010",
				"100110101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100010101010",
				"100010011010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100111",
				"010001100111",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"010001010110",
				"010001010110",
				"010001010110",
				"010001010110",
				"010001010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001000110011",
				"001000110010",
				"001000110010",
				"001000110011",
				"001100110011",
				"001101000011",
				"010001000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001000100",
				"010001000100",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"001101000011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000011",
				"010001000100",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000011",
				"010001000100",
				"010101010100",
				"010001000100",
				"010000110011",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001101010101",
				"011010001000",
				"100110101011",
				"101010111100",
				"101111001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101000100",
				"001101010101",
				"001101010100",
				"001101000100",
				"001001000100",
				"001001000011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000110011",
				"001101000011",
				"001101000100",
				"010001000100",
				"010001010100",
				"001101000100",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"001101000011",
				"001101000011",
				"010001000100",
				"001101000011",
				"001101000011",
				"010001000011",
				"001100110011",
				"001100110010",
				"001100110011",
				"010001000100",
				"010101000100",
				"010000110011",
				"010000110011",
				"010001000011",
				"010101000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"001100110011",
				"001100110010",
				"010001000011",
				"010001000100",
				"010001000100",
				"001101000011",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001000100010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100100010",
				"001100110010",
				"001100100010",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100110011",
				"010101100111",
				"100010101010",
				"100110111011",
				"101110111100",
				"101111001100",
				"110011001101",
				"110011001100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101001",
				"100110101001",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101111000",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101010110",
				"001101010110",
				"010001010101",
				"010001100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101010101",
				"001101010101",
				"001101010100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000011",
				"001000110011",
				"001000110011",
				"001001000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"010001010100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001101000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001100110010",
				"001000100010",
				"001100100010",
				"010000110011",
				"010101000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000011",
				"001101000011",
				"001101000011",
				"001100110010",
				"001000110010",
				"001000110010",
				"001100110011",
				"001100110011",
				"001101000011",
				"010001000011",
				"010001000100",
				"001100110010",
				"001000100001",
				"001000100001",
				"001100110010",
				"010001000011",
				"010101000100",
				"010101010100",
				"010001000011",
				"010001000011",
				"001100110011",
				"001100110010",
				"001100110010",
				"001000100001",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001101000100",
				"011010001000",
				"100110101010",
				"101010101011",
				"101110111100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010011010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"001101111000",
				"001101110111",
				"001101110111",
				"001101111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101010100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"010001010100",
				"010001010100",
				"001101000100",
				"001101000011",
				"001101000011",
				"001101000100",
				"010001000100",
				"010001000100",
				"001101000100",
				"001101000011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000011",
				"010001000011",
				"010001000011",
				"001100110011",
				"001100110010",
				"001100110010",
				"001100110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001010100",
				"010001010100",
				"001101000011",
				"001000110010",
				"001100110011",
				"001101000011",
				"001101000100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101000100",
				"001100110011",
				"001100110011",
				"010001000011",
				"010101000100",
				"010101000100",
				"010101000100",
				"010101000100",
				"010001000011",
				"010001000011",
				"001100110010",
				"001100100010",
				"001100110011",
				"001100110011",
				"001100110010",
				"001100100010",
				"001000100010",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"010001010110",
				"100010011001",
				"100110101010",
				"101010111100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"001101111000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"001101111000",
				"001101111000",
				"001101111000",
				"010001111000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101000100",
				"001001000011",
				"001001000011",
				"001000110011",
				"001101000100",
				"001101010100",
				"010001010101",
				"010001010100",
				"001101000011",
				"001000110010",
				"001001000011",
				"010001010100",
				"010001010100",
				"001101000100",
				"001101000011",
				"001101000011",
				"010001000011",
				"010001000100",
				"010001000011",
				"001101000011",
				"010001000011",
				"001100110011",
				"001100110011",
				"010001000011",
				"010001000011",
				"010001000100",
				"010001000011",
				"001100110011",
				"010001010100",
				"010101010101",
				"010001010100",
				"001101000011",
				"001100110011",
				"001101000011",
				"010001010100",
				"010001010100",
				"010101100101",
				"010101100101",
				"010101010101",
				"010101010100",
				"010001010100",
				"010001000100",
				"001100110011",
				"001000100010",
				"001100110011",
				"010001000011",
				"010101010101",
				"011001100101",
				"010101010101",
				"010101000100",
				"010101000100",
				"010001000011",
				"001000010001",
				"000100000000",
				"000100010000",
				"001100100010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001100110010",
				"001000010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000110011",
				"011001110111",
				"100010011010",
				"101010111011",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010001111000",
				"001101111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"001101111000",
				"001101111000",
				"001101111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000101",
				"001101000101",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001000110011",
				"001001000100",
				"001101000100",
				"001101010100",
				"001101010101",
				"001101010101",
				"001101000100",
				"001001000011",
				"001001000011",
				"001101000100",
				"001101010100",
				"010001010101",
				"010001010100",
				"001001000011",
				"001000110010",
				"001001000011",
				"001101010100",
				"010001010100",
				"001101000100",
				"001101000011",
				"001101000011",
				"010001000100",
				"010001000100",
				"001100110011",
				"001100110010",
				"001100110010",
				"001100110010",
				"010000110011",
				"010101010100",
				"010101010101",
				"010001000100",
				"010001000011",
				"010001000011",
				"010101010101",
				"010101010101",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010100",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110010",
				"001000110010",
				"010001000100",
				"010001000100",
				"010101000100",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101000100",
				"010001000100",
				"001000010001",
				"000100000000",
				"000100010001",
				"001100100010",
				"001100110010",
				"001100110011",
				"010000110011",
				"010001000011",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"010001010101",
				"011110001000",
				"100110101010",
				"101010111100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110011010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"001101111000",
				"001101111000",
				"001101111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001001000100",
				"001001000100",
				"001000110100",
				"001000110100",
				"001001000100",
				"001001000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"001101010100",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101010100",
				"010001010101",
				"010001010101",
				"001101010100",
				"001001000011",
				"001000110010",
				"001001000011",
				"001101010100",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001010100",
				"010001010100",
				"010001000011",
				"001100110011",
				"001100100010",
				"001100100010",
				"001100110010",
				"010101010100",
				"011001100101",
				"011001100101",
				"010001010100",
				"010001010100",
				"010101010101",
				"011001100101",
				"010001000100",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010101100101",
				"010101100101",
				"010001010101",
				"001001000011",
				"000100110010",
				"001000110011",
				"001101010100",
				"010001100101",
				"010101100110",
				"010101010101",
				"010101010101",
				"010101010100",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010100",
				"010000110011",
				"001100110011",
				"010000110011",
				"010001000011",
				"010001000011",
				"010001000100",
				"010101010100",
				"010101010100",
				"010001010100",
				"001100110011",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"010101100110",
				"100010011001",
				"101010111011",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"001101111000",
				"001101111000",
				"001101111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101010110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001001000100",
				"001001000100",
				"000100110100",
				"000100110011",
				"001001000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001000100",
				"001101000100",
				"001101000100",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101000100",
				"001000110011",
				"001001000011",
				"001101000100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000011",
				"010000110011",
				"010000110011",
				"010101000100",
				"011001100101",
				"011101110110",
				"011001100110",
				"010101100101",
				"010101100101",
				"011001100110",
				"011001010101",
				"010000110011",
				"001000100010",
				"001100110010",
				"010001000100",
				"010001000100",
				"010001010100",
				"010001010101",
				"010101100101",
				"010101100110",
				"010001100101",
				"001001000011",
				"000100110011",
				"001001000011",
				"010001100101",
				"010101100110",
				"010101100101",
				"010101010101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010001000100",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010100",
				"010001010100",
				"010101010101",
				"010001000100",
				"010001000100",
				"010001000011",
				"001000100010",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001101000100",
				"011101111000",
				"100110101010",
				"101010111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110011010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"001101111000",
				"001101111000",
				"001101111000",
				"001101111000",
				"001110001000",
				"010010001000",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001001000101",
				"001001000100",
				"001001000100",
				"001001000101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001001000100",
				"001001000100",
				"001001000100",
				"001101010101",
				"010001010101",
				"010001100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"001101000011",
				"001000110011",
				"001101000100",
				"010001010100",
				"010101100101",
				"010001010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010100",
				"010101010100",
				"010101000100",
				"010101000100",
				"010101000100",
				"011001010101",
				"011101110110",
				"011101110111",
				"011101110110",
				"011001110110",
				"010101100101",
				"010101100101",
				"010001010101",
				"001100110011",
				"001000110011",
				"010001010101",
				"011001100110",
				"010101010101",
				"010101010101",
				"010101100110",
				"010001010101",
				"010101100110",
				"010101100110",
				"001101010100",
				"001101000100",
				"001101010100",
				"010001010101",
				"010001100101",
				"010101100110",
				"010001010101",
				"010001010101",
				"010101100110",
				"011001100110",
				"011001100110",
				"010001010100",
				"001100110011",
				"001100110011",
				"001101000011",
				"010001000100",
				"010101010100",
				"010101100101",
				"010101100101",
				"010101100101",
				"010001010100",
				"010001010100",
				"010001000100",
				"010001000011",
				"001100110011",
				"001000100001",
				"000100010001",
				"000100010001",
				"001000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"010001010101",
				"011110011001",
				"100110101011",
				"101010111011",
				"101010111100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"001101111000",
				"001101111000",
				"001101111000",
				"001101111000",
				"010010001000",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"001101010110",
				"001101010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001001000101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010101100110",
				"010001010101",
				"001101000100",
				"001001000100",
				"001001000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001000100",
				"010001010100",
				"010101100101",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010101010101",
				"010101010100",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"010001010101",
				"001101000100",
				"001101000100",
				"010001100110",
				"010001100110",
				"011001110111",
				"011010000111",
				"010101110110",
				"011001110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101010101",
				"001101000100",
				"010101010101",
				"011001100110",
				"010101010110",
				"010101100110",
				"010101100110",
				"011010000111",
				"011001110111",
				"010001010101",
				"010001000100",
				"010001010101",
				"001100110011",
				"001000110010",
				"001000110011",
				"001101000011",
				"010001010100",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010001010100",
				"010001000100",
				"001101000011",
				"001000100010",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110010",
				"001000100010",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000100011",
				"010101100110",
				"011110001000",
				"100110101010",
				"101010111011",
				"101110111011",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010101100101",
				"010101100110",
				"010001010101",
				"010001010101",
				"010101010101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101110110",
				"010101100101",
				"010101010101",
				"010001010100",
				"010101010100",
				"010001000100",
				"011001100101",
				"010001000100",
				"010101100101",
				"011001100110",
				"010101100101",
				"010001010100",
				"001101010100",
				"010101100101",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"011101110111",
				"010101100110",
				"010001000100",
				"001100110011",
				"010101010101",
				"011101100111",
				"011001100110",
				"011001100111",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001010101",
				"001000110011",
				"001101000100",
				"010001010101",
				"010101010101",
				"010101100101",
				"010001100101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010101",
				"010101100101",
				"010101100110",
				"010101010101",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001010100",
				"010101010101",
				"010101010100",
				"010001000100",
				"001100110011",
				"001000110010",
				"000100100001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"010001010101",
				"011110001000",
				"100010011010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100110",
				"001101010101",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100110",
				"001101010101",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010101010101",
				"011001100110",
				"010101100110",
				"010001010101",
				"010001000100",
				"010001010101",
				"010101100101",
				"010101100110",
				"011001110110",
				"011001100110",
				"010101010101",
				"010001000100",
				"010001000100",
				"010101010101",
				"011001100110",
				"010001010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"010101100101",
				"010001010101",
				"010001100101",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"010101100110",
				"010001010101",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"011001100110",
				"011001100111",
				"011001100110",
				"011001110111",
				"010101110110",
				"010001100110",
				"010101110110",
				"010101110111",
				"011001110111",
				"010001010101",
				"001000110011",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101010101",
				"010001000100",
				"001101000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010001010101",
				"010001000100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000100011",
				"010101100110",
				"011110001000",
				"100110101010",
				"101010101011",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110111",
				"010001100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101100101",
				"010001000100",
				"010001000100",
				"010101100101",
				"011001110110",
				"010101100110",
				"010101100110",
				"011001110110",
				"010101100110",
				"010001010100",
				"010001010100",
				"011001100110",
				"010101100101",
				"010001000100",
				"001101000100",
				"010001010100",
				"010101100110",
				"011010000111",
				"010101110110",
				"010001010101",
				"010101100110",
				"010101110111",
				"011001111000",
				"010101100110",
				"010001100110",
				"010001010110",
				"010001010101",
				"010101100111",
				"011001100111",
				"010101100111",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010001100110",
				"010101110110",
				"011001110111",
				"011001110111",
				"010001010101",
				"001000110011",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100101",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101100110",
				"010101100101",
				"011001110111",
				"011001100110",
				"010001010101",
				"001000100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001100110100",
				"010101100110",
				"100010011001",
				"100110101010",
				"101010101011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110011010",
				"011110011001",
				"011110011001",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"001110001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100101",
				"010001100110",
				"010101110110",
				"011001110111",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010101",
				"010101100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"010101100110",
				"010101100110",
				"011001110110",
				"001101000100",
				"001000110011",
				"001101010100",
				"010101110110",
				"011001110111",
				"011001110111",
				"010101110111",
				"011001110111",
				"011110001000",
				"011101111000",
				"011001110111",
				"010101010110",
				"010101010110",
				"011001110111",
				"011001110111",
				"100010011001",
				"011110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010110000111",
				"010110001000",
				"010010000111",
				"010001110110",
				"010001110110",
				"010001100110",
				"010101110110",
				"010101110110",
				"011001110111",
				"010101110110",
				"010001010101",
				"010101100110",
				"011001100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100101",
				"010101110110",
				"010001100110",
				"010101100110",
				"010101110110",
				"010001010101",
				"001000110011",
				"001000110011",
				"001100110011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001001000011",
				"001001000011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001000110011",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000010001",
				"000100010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001101000100",
				"011001110111",
				"100010011001",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"001101100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"001101010101",
				"010001100101",
				"010101110110",
				"010101110111",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010001010101",
				"010101100110",
				"011001100110",
				"011001100110",
				"011001110110",
				"011010000111",
				"011001110111",
				"010001100101",
				"001000110011",
				"001001000100",
				"010101100110",
				"011001110111",
				"011010000111",
				"011010001000",
				"011010000111",
				"011001110111",
				"100010011001",
				"011101110111",
				"010101010110",
				"011001100110",
				"100010001001",
				"100110101010",
				"100010011001",
				"011110001000",
				"010101110111",
				"010001110111",
				"010110000111",
				"010110000111",
				"010010000111",
				"010110011000",
				"010110011001",
				"010110011000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"011001110111",
				"011001110111",
				"010101010101",
				"010101100110",
				"011001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101000100",
				"001000110011",
				"001000110011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101010100",
				"001101010100",
				"001101010100",
				"001101000100",
				"001001000100",
				"001001000011",
				"001000110011",
				"000100100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"001100110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"010001000101",
				"011101111000",
				"100110011010",
				"101010101011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101010",
				"100010101010",
				"100010101010",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101100111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010001100110",
				"001101100101",
				"010001100110",
				"010101110110",
				"010101110111",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001100110",
				"010101110110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010101100110",
				"011001110110",
				"011001100110",
				"011001110111",
				"011010000111",
				"010101110110",
				"010001010101",
				"001101010100",
				"010001100110",
				"011010000111",
				"010101110111",
				"010101110111",
				"011110001000",
				"011001111000",
				"010001010110",
				"010101100110",
				"011001110111",
				"011101111000",
				"011110001001",
				"100010011001",
				"011110001001",
				"011010001000",
				"011010001000",
				"010001100110",
				"010001100110",
				"010110001000",
				"010110001000",
				"010010000111",
				"010010000111",
				"010010001000",
				"010110001000",
				"011010011000",
				"011010001000",
				"011010001000",
				"011001110111",
				"011001110111",
				"010001010101",
				"001101000100",
				"010001010101",
				"011001100110",
				"011001110111",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001000100",
				"010001000100",
				"010001010101",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"001101000011",
				"001100110011",
				"001000100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000000000",
				"000000000001",
				"001000100011",
				"010101100110",
				"100010001001",
				"100110101010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101010",
				"100010101010",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010101111000",
				"010101111000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110000111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010101110111",
				"011010000111",
				"010101110110",
				"010001010101",
				"001101010101",
				"010101100110",
				"010101110110",
				"010001100101",
				"010001100101",
				"010101100101",
				"010101100110",
				"010101100110",
				"011001100110",
				"011001110111",
				"011001110111",
				"010101110110",
				"010001100101",
				"010001010101",
				"010101110110",
				"010101110111",
				"011010001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001010101",
				"010001100110",
				"011010001000",
				"011010001000",
				"011110001001",
				"011010001000",
				"010001110111",
				"011010001000",
				"011010011001",
				"010001110111",
				"001101100101",
				"010001110111",
				"010110001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110000111",
				"011001110111",
				"011001110110",
				"011001110111",
				"011110001000",
				"011110001000",
				"010101010110",
				"010001000100",
				"011001100111",
				"011110001000",
				"011110001001",
				"011110001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101100110",
				"010001010101",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010001100110",
				"010001100101",
				"010001100101",
				"001101100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010101100101",
				"010101100101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010101010101",
				"010001010101",
				"010001000100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110011",
				"011001100111",
				"100010001001",
				"100110101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"110010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101110101011",
				"101110111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"101010101011",
				"101010101011",
				"100110101011",
				"100110101010",
				"100110101011",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100110",
				"001101100111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110000111",
				"010001110111",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001110110",
				"011010000111",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100101",
				"010101100110",
				"011001110111",
				"010101100110",
				"010001010101",
				"010001100101",
				"010101100110",
				"011001100110",
				"010001000100",
				"010101110110",
				"011010000111",
				"010101100110",
				"010101100110",
				"010101100101",
				"011001110111",
				"011010000111",
				"010110011000",
				"010110011000",
				"010110001000",
				"011110011001",
				"011110001001",
				"010001010110",
				"010001010101",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"001101100110",
				"010001110111",
				"011010001000",
				"010101110111",
				"011001111000",
				"011101111000",
				"011001100111",
				"011101110111",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100111",
				"011001100111",
				"011001111000",
				"011010001000",
				"010101111000",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010001110111",
				"010110001000",
				"010101110111",
				"010001110111",
				"011010001000",
				"011110011001",
				"010101110111",
				"001101100110",
				"001101100110",
				"010001110111",
				"001001100101",
				"010110000111",
				"010110000111",
				"010001110110",
				"010101110111",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"001101010101",
				"001101000100",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110111",
				"011001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110111",
				"011001110111",
				"011001100110",
				"010001010101",
				"001100110011",
				"001000100010",
				"001000100010",
				"001100100010",
				"001100100010",
				"001000010001",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001101000100",
				"011001100111",
				"100010001001",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"110010111010",
				"110010111010",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101010",
				"100110101011",
				"100110101010",
				"100110101010",
				"100110101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"011010000111",
				"010110000111",
				"010101110110",
				"010001100110",
				"010101100110",
				"010101110111",
				"011001110110",
				"010101100110",
				"010001100101",
				"010101100101",
				"010101100101",
				"011001100101",
				"010101010101",
				"010101100110",
				"010101110110",
				"010101100110",
				"010101100101",
				"010101100110",
				"011010000111",
				"011010011000",
				"011010011000",
				"011010011001",
				"011010011001",
				"011110011001",
				"011010001000",
				"010001010110",
				"010101100110",
				"011010001000",
				"010110001000",
				"010101111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011110011001",
				"011110001001",
				"011001100111",
				"011101101000",
				"100110001001",
				"100110011001",
				"100010000111",
				"011101110111",
				"011101111000",
				"100010001000",
				"100010001001",
				"011110001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010001110111",
				"001101100110",
				"010001110110",
				"001101110110",
				"010001110110",
				"010001100110",
				"010001110110",
				"011010000111",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010001100110",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001010101",
				"010101010101",
				"010001010101",
				"010101010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101010101",
				"010101010101",
				"010101010100",
				"010101010100",
				"010101010100",
				"010001000100",
				"010000110011",
				"001100100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001101000100",
				"011001100111",
				"100010011001",
				"100110101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"110010111010",
				"110010111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110101011",
				"101110101011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"100110101010",
				"100110101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010110001000",
				"010101110111",
				"010001110110",
				"010001100110",
				"010101110111",
				"010110000111",
				"011010000111",
				"010101110111",
				"010001100110",
				"010001100110",
				"011001110111",
				"011010000111",
				"011001110110",
				"010101110110",
				"010101100110",
				"010101100101",
				"010101010101",
				"010101010101",
				"011001100110",
				"010101010101",
				"010101010101",
				"011001100110",
				"010001010101",
				"010101100110",
				"011010011000",
				"010110000111",
				"011010011000",
				"011110011001",
				"011010001000",
				"011001111000",
				"010101110111",
				"010101100111",
				"011010001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110001000",
				"011001111000",
				"011001110111",
				"011101111000",
				"100010001001",
				"100110001010",
				"101010101011",
				"101010111011",
				"100110111010",
				"100110111011",
				"100110101010",
				"100010011001",
				"011110001001",
				"011010001000",
				"010110001000",
				"011010011001",
				"010110001001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"011010001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"011010011001",
				"011110011001",
				"011010001000",
				"010001100110",
				"010101110111",
				"011110011001",
				"011010001000",
				"010101110110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110111",
				"010101100110",
				"010001010101",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001000101",
				"001101000100",
				"001101010100",
				"001001000100",
				"001001000011",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010100",
				"001101000011",
				"000100100001",
				"001000100010",
				"001000110010",
				"001101000011",
				"010001000100",
				"010001010101",
				"010001000100",
				"001100110011",
				"000100010001",
				"000100010001",
				"000100010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100010",
				"001101000100",
				"010101100110",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010101011",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101010",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111011",
				"100110111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010111011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011010011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010101010",
				"011110101010",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010101110111",
				"010110000111",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100101",
				"010101100110",
				"011010000111",
				"011010000111",
				"011001110110",
				"011001110111",
				"011001110110",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010001000100",
				"011001100101",
				"011001110110",
				"010001010100",
				"010001110110",
				"011010011000",
				"011010001000",
				"011110001000",
				"011001111000",
				"010101100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010011001",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011001111000",
				"011001110111",
				"011101111000",
				"011001100111",
				"010101100110",
				"011001110111",
				"100010011010",
				"100110101011",
				"100110101011",
				"100010011010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010001001",
				"010110001001",
				"010001111000",
				"010001111000",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010101010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010001110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010001010101",
				"010101010110",
				"010101010101",
				"010001010101",
				"010001000100",
				"001101000100",
				"001001000100",
				"001101010100",
				"001101010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110111",
				"010101110111",
				"010001010101",
				"001101000100",
				"010001010101",
				"010001100110",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010101100101",
				"010001100101",
				"010001010100",
				"010001010101",
				"010001010100",
				"001101000100",
				"001101000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001000110011",
				"001101000011",
				"001100110011",
				"001000110010",
				"000100100001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110011",
				"010101010101",
				"011101110111",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"100110101011",
				"101010101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011010011010",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"011010000111",
				"011001110111",
				"011001110110",
				"011110000111",
				"011001110111",
				"011001100110",
				"011001100110",
				"010101110110",
				"001101000011",
				"010000110011",
				"011101100110",
				"011101110111",
				"001101010100",
				"010001110110",
				"011010011000",
				"011110011001",
				"011101111000",
				"010101100110",
				"010101100111",
				"011110011001",
				"011110101010",
				"011010011001",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"100010011001",
				"100010001001",
				"010101010110",
				"011001010110",
				"100010001001",
				"100110101011",
				"011110101010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011010",
				"010010001001",
				"001110001000",
				"010010001000",
				"010010011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010110011001",
				"011010011001",
				"010110001000",
				"010010011001",
				"010010011000",
				"010110101010",
				"011010101010",
				"010110001000",
				"010001110111",
				"011010001000",
				"011110001001",
				"010001000101",
				"001000010010",
				"001100100011",
				"010101000101",
				"010101010101",
				"010101100110",
				"010101100110",
				"010101110111",
				"010101110111",
				"011001110111",
				"010101110111",
				"010101100110",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010001110110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"001101100101",
				"010001100101",
				"010001100101",
				"010101100110",
				"010101110110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001010101",
				"001101010100",
				"001101000011",
				"001000110011",
				"001000110010",
				"001000100010",
				"000100100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000100010",
				"001101000100",
				"011001100110",
				"100010001000",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101011",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"011010000111",
				"011001110111",
				"010101110110",
				"011001110110",
				"011001110111",
				"011001110110",
				"011001110110",
				"011001110110",
				"010101100101",
				"001000110010",
				"010001000100",
				"011101110111",
				"011110001000",
				"010001100101",
				"011010000111",
				"011110011001",
				"010101100110",
				"010101010110",
				"010101100110",
				"011110001001",
				"011110101010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011110011001",
				"011110011001",
				"100010011001",
				"011101111000",
				"010101010110",
				"011001100111",
				"100010001001",
				"011010001001",
				"010110001000",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110101010",
				"010010011001",
				"010010001001",
				"001110001000",
				"010010011001",
				"010110011010",
				"010110011001",
				"010110001001",
				"011010011010",
				"011010011001",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010011000",
				"010110001000",
				"010110001000",
				"011110001001",
				"100010011001",
				"100110001001",
				"010101000110",
				"001000010011",
				"010101000110",
				"011101111000",
				"011101111000",
				"011110001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"010010000111",
				"001101110110",
				"001101100110",
				"001101110110",
				"010010000111",
				"010001110111",
				"001101100110",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110110",
				"010001110110",
				"010001110110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100101",
				"010101100101",
				"010101010101",
				"010001010100",
				"001101000011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110011",
				"010101010101",
				"011101110111",
				"100010011001",
				"100110011010",
				"101010101010",
				"101010101011",
				"101010101010",
				"101010101011",
				"101010111011",
				"101110111011",
				"101110101011",
				"101110101011",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"100010111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110110",
				"011001110111",
				"011001110110",
				"011001110110",
				"011001110110",
				"011101110111",
				"011110000111",
				"010001010100",
				"001001000011",
				"010101100101",
				"011110000111",
				"100010011000",
				"010101100110",
				"010101100110",
				"011001110111",
				"001101000100",
				"010101010110",
				"011001111000",
				"011110101010",
				"011010011001",
				"010001110111",
				"010110001001",
				"011010011001",
				"010110011001",
				"010110101001",
				"011010101001",
				"011010011001",
				"011110011001",
				"011110001000",
				"011101111000",
				"011101111000",
				"010101010110",
				"010101110111",
				"011110011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010010011001",
				"001110001000",
				"010001111000",
				"010001111000",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"001101111000",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"011101111000",
				"011101111000",
				"011001100111",
				"010001000101",
				"001100110100",
				"001101000100",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010001111000",
				"010001111000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110011001",
				"010110011000",
				"010110011001",
				"010010001000",
				"001101100110",
				"001101100110",
				"010001110111",
				"010110000111",
				"010110000111",
				"011010000111",
				"011010000111",
				"011010000111",
				"010110000111",
				"010101110111",
				"010101110110",
				"010001100101",
				"010101110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100101",
				"010001010100",
				"001100110011",
				"001000100010",
				"000100010001",
				"000000000000",
				"000100000000",
				"000100000000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000100011",
				"010001010101",
				"011001110111",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110011011",
				"010010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010010000111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"011001110111",
				"011001110111",
				"010101100110",
				"011001100110",
				"011110000111",
				"011110000111",
				"001101000011",
				"010001010100",
				"011110000111",
				"011001110111",
				"011110001000",
				"010101010101",
				"001100110100",
				"001100110100",
				"010101010110",
				"011001111000",
				"011110011001",
				"011010101010",
				"010110001000",
				"010010001000",
				"011010011001",
				"011010011001",
				"011010101001",
				"011010101001",
				"011110011001",
				"011110011001",
				"011110001000",
				"011101110111",
				"011001100111",
				"011001010110",
				"100010011001",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010110001001",
				"010110011010",
				"010110011010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011110011001",
				"011001111000",
				"010101100111",
				"010101010110",
				"010000110101",
				"001100100100",
				"001000100011",
				"010101100110",
				"011010001000",
				"010110001000",
				"010010001000",
				"010010011000",
				"010010011001",
				"010010011000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010010001000",
				"010110011000",
				"011010101001",
				"011010011001",
				"010001110111",
				"001101100110",
				"010001110111",
				"010001110111",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110111",
				"011010000111",
				"011010000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001010101",
				"010001010100",
				"001000100010",
				"001000100010",
				"001000110010",
				"001000110010",
				"001000100010",
				"001000100010",
				"001000100001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"010001000100",
				"011001110111",
				"100010001001",
				"100010011001",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110101011",
				"100010111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"010110101011",
				"010110101011",
				"010010011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"011010011000",
				"010101110111",
				"010001110110",
				"011010000111",
				"011010000111",
				"011001110110",
				"010101100110",
				"011001110110",
				"011101110111",
				"011001110110",
				"010001100101",
				"010001100101",
				"011110011000",
				"010101110110",
				"100010011000",
				"010001000101",
				"000000000001",
				"010001000101",
				"011110001000",
				"011110011010",
				"011010011001",
				"011010011001",
				"011110101011",
				"010110001000",
				"011110011001",
				"100110111011",
				"100010101010",
				"011110011001",
				"011001110111",
				"011001100111",
				"011101010111",
				"011001010110",
				"011101100111",
				"100110001001",
				"100110101011",
				"100010101011",
				"011010011010",
				"010110011001",
				"011010011010",
				"010110011010",
				"010110001001",
				"011110011010",
				"011110011010",
				"011010001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110001001",
				"011001111000",
				"100110101011",
				"011110001001",
				"011110011010",
				"011010001000",
				"010101110111",
				"010101100111",
				"010001010110",
				"010001010110",
				"010001000101",
				"010001000101",
				"010001000101",
				"010101010110",
				"010101100111",
				"011010011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110101001",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011110011001",
				"011110011001",
				"010101110111",
				"001101100110",
				"010101110111",
				"011001110111",
				"011001110111",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101010100",
				"010001010101",
				"001101010100",
				"001101010100",
				"001101000100",
				"001101010100",
				"010001010101",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000000010000",
				"000100010001",
				"000100100001",
				"001000100010",
				"000100010001",
				"000000010000",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000100010",
				"010001010101",
				"011001100111",
				"100010011001",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101010101010",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110101010",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010110001000",
				"011010011000",
				"011010001000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101110110",
				"010101100110",
				"011001110111",
				"011110000111",
				"011110001000",
				"011010000111",
				"011010000111",
				"011110011000",
				"011110001000",
				"100010001000",
				"001100100011",
				"001000010010",
				"011001100111",
				"011010001001",
				"011010101010",
				"011010101010",
				"011010101010",
				"100010111011",
				"011010011001",
				"011110011001",
				"100010011010",
				"011101111000",
				"011001100111",
				"010101010110",
				"011001100111",
				"100010001001",
				"100010001001",
				"100010001001",
				"100010011010",
				"100110101011",
				"011110011010",
				"011010011001",
				"011010011010",
				"011010011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011110101010",
				"011110101011",
				"011010101010",
				"010110011001",
				"010110001000",
				"010101111000",
				"010101111000",
				"011110001000",
				"011101111000",
				"010001000101",
				"011001100111",
				"010101100111",
				"010101010110",
				"010001000101",
				"010001010110",
				"010001010110",
				"010001100111",
				"010101110111",
				"011001111000",
				"011010001000",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101110111",
				"011010001000",
				"011110011001",
				"011110001001",
				"011001111000",
				"010101110111",
				"011110001000",
				"011110001000",
				"011110001000",
				"011001110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001010101",
				"001101000101",
				"001001000100",
				"001101000101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010100",
				"001101010100",
				"001101010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001000011",
				"001101000100",
				"001101000011",
				"001000110011",
				"001000110011",
				"001000110011",
				"000100110010",
				"000100100010",
				"000100100010",
				"001000110010",
				"001000110010",
				"001000110011",
				"001000110011",
				"000100100010",
				"000100010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"001101000100",
				"011001110111",
				"011110001000",
				"100110011001",
				"100110101010",
				"101010101011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101110111",
				"011010000111",
				"011010001000",
				"011010001000",
				"010101110110",
				"010101110110",
				"011001110111",
				"100010011000",
				"100110101001",
				"100010101001",
				"011110011000",
				"011110011000",
				"100010011001",
				"100001111000",
				"001000010010",
				"001100110100",
				"011001111000",
				"011010011001",
				"010110101001",
				"011010101010",
				"011010011001",
				"011110101010",
				"011110011001",
				"011001111000",
				"010101100111",
				"011001010110",
				"011101010111",
				"011101100111",
				"011110001000",
				"100010011010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010101011",
				"011010001001",
				"011010001001",
				"011110011010",
				"011010001001",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110101010",
				"011010111011",
				"011110111010",
				"011010011001",
				"011010001000",
				"011001110111",
				"011110001001",
				"001100110100",
				"001100110100",
				"010001000101",
				"010101100111",
				"010101100111",
				"011001111000",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110001001",
				"010001111000",
				"010110001001",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101110111",
				"010001100111",
				"011001111000",
				"011110011001",
				"011010001000",
				"010001010101",
				"011001100111",
				"011001110111",
				"011110001000",
				"011110001000",
				"011010001000",
				"011001111000",
				"011001111000",
				"010101111000",
				"010101111000",
				"010101110111",
				"010101111000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001010110",
				"010001010110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"001101010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"001101000011",
				"001000110011",
				"000100100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001101000100",
				"010101100110",
				"100010001000",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110101011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010111011",
				"100110111011",
				"100110111011",
				"100010101011",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111100",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010101010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010011001",
				"011110101001",
				"011010011001",
				"010110001000",
				"010101110111",
				"011010001000",
				"011010011000",
				"011010001000",
				"011001110111",
				"011010000111",
				"011110001000",
				"100010011001",
				"100110111010",
				"011110101001",
				"011110101001",
				"100010011001",
				"100010001001",
				"011001010110",
				"001000010010",
				"010101010110",
				"011010001000",
				"011010101010",
				"010010101001",
				"011010101010",
				"010110011001",
				"011110001001",
				"011110001001",
				"010001010110",
				"001100110100",
				"011101100111",
				"100101111001",
				"100110011010",
				"100010011010",
				"011110101010",
				"011010011010",
				"011010101010",
				"011110111011",
				"011110101010",
				"011010001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010101010",
				"010010101010",
				"010010101001",
				"010110101001",
				"010110011001",
				"011010011001",
				"011110011001",
				"100010101010",
				"100010011010",
				"001100110100",
				"001101000100",
				"010101100111",
				"011110001001",
				"011110011001",
				"011010001001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001000",
				"010010011001",
				"010010011001",
				"010110001001",
				"011010101010",
				"011010011001",
				"010101111000",
				"010110001000",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011110101010",
				"011110101010",
				"011110011001",
				"010101111000",
				"010001100110",
				"010101110111",
				"011110001000",
				"011001111000",
				"011001111000",
				"011110001000",
				"100010011001",
				"011110011001",
				"011110001001",
				"011010001001",
				"011010001001",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001001",
				"011010001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001001",
				"011010001000",
				"010101111000",
				"010101110111",
				"010101110111",
				"011010001000",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110111",
				"010101110110",
				"010101110111",
				"010101110110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101100110",
				"011001100110",
				"010101100110",
				"010101010101",
				"010001010100",
				"001101000100",
				"001000110011",
				"000100100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001100110011",
				"010101100110",
				"011110001000",
				"100110011001",
				"100110101010",
				"101010111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110101011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010010011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110011000",
				"010110011000",
				"011010011000",
				"011110101001",
				"011110101001",
				"011010011000",
				"010110001000",
				"010110000111",
				"011010011000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011110001000",
				"011110001000",
				"011110011001",
				"100010101010",
				"011010000111",
				"100010101001",
				"100110101010",
				"011101110111",
				"010001000100",
				"010001000100",
				"011010001000",
				"011010011001",
				"010110101010",
				"010010011001",
				"011010101010",
				"011010011001",
				"011110011001",
				"100010011010",
				"010101010110",
				"001101000100",
				"011110001001",
				"100010011010",
				"100010011010",
				"011110011010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010010101010",
				"010010101010",
				"010110101010",
				"010110101001",
				"010110101001",
				"011010011001",
				"011110101010",
				"100010011010",
				"010101100110",
				"001000110011",
				"010101100111",
				"011110011010",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010001111000",
				"001101111000",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"010110001000",
				"010101110111",
				"011001111000",
				"011001110111",
				"011001110111",
				"011010001000",
				"011110001001",
				"011010001001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101110111",
				"010110001000",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010001110111",
				"010001100110",
				"010001110111",
				"010101111000",
				"010101110111",
				"010101110111",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001110110",
				"010101110111",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001010101",
				"010001000100",
				"001101000100",
				"010001000100",
				"001101000100",
				"001100110011",
				"001100110011",
				"001000110011",
				"001000110010",
				"001000110010",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110011",
				"010101010101",
				"011101110111",
				"100010011001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"110010111100",
				"110010111100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011000",
				"011010011000",
				"011010011001",
				"011010101001",
				"011010011000",
				"010110001000",
				"010110000111",
				"010110001000",
				"011110011001",
				"011010011000",
				"011010011000",
				"011110011001",
				"011110001000",
				"011110001000",
				"011110011001",
				"011110011000",
				"011110001000",
				"100010011001",
				"100010001000",
				"010101010101",
				"010001010101",
				"011001111000",
				"011110101010",
				"011010011010",
				"011010101010",
				"010110101010",
				"011010101010",
				"011010101001",
				"011110011001",
				"100010011010",
				"010101010110",
				"010001010101",
				"011110001001",
				"011110011010",
				"011110101010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010111011",
				"010010011001",
				"010010011001",
				"010110101010",
				"011010101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"011010101010",
				"011110101010",
				"011110101010",
				"011010001000",
				"011001111000",
				"010001010101",
				"001100110100",
				"010001010110",
				"100010011010",
				"011110011010",
				"010110011001",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101100110",
				"010101100110",
				"010101100111",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010001110111",
				"010001100111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110000111",
				"011010001000",
				"011010001000",
				"010110000111",
				"011010000111",
				"011010000111",
				"011010000111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"011001110110",
				"010101100101",
				"010001000100",
				"001100110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000100010",
				"010001000100",
				"011001100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110101010",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100010101010",
				"100010101010",
				"011110101010",
				"011110101010",
				"011110101011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101011",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011000",
				"011010011001",
				"011010101001",
				"011010011001",
				"010110001000",
				"010001110111",
				"010110000111",
				"011010011001",
				"011110101001",
				"011010011000",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110001000",
				"100010011001",
				"100010001001",
				"011001100111",
				"010001010101",
				"010101110111",
				"011110101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"100010011001",
				"010101010110",
				"010101010110",
				"011110011010",
				"011110101011",
				"011110101011",
				"011110011010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110011011",
				"100010011011",
				"100010011011",
				"100010011011",
				"011110011010",
				"011001111000",
				"010001010110",
				"010001000101",
				"010001000101",
				"010001000101",
				"011001010110",
				"100110011010",
				"100110101011",
				"011010001001",
				"010110011010",
				"010110101010",
				"010010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"010110001001",
				"001101100111",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011001",
				"011110011001",
				"011001110111",
				"010001010101",
				"001101000100",
				"010101010110",
				"011110001000",
				"011110001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010101110111",
				"010001100110",
				"001101010101",
				"001001000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000011",
				"001101000100",
				"001101000100",
				"010001010101",
				"010101010101",
				"010101100101",
				"010101010101",
				"010001010100",
				"001100110011",
				"001000100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"001100110100",
				"010101010101",
				"011001110111",
				"011101111000",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101110111100",
				"101110111100",
				"101010111100",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110101010",
				"100010101010",
				"100010101010",
				"100010101011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"100010111011",
				"100010111011",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010101001",
				"011110101001",
				"011010011001",
				"010110000111",
				"010001110111",
				"010110011000",
				"011110101001",
				"011110101001",
				"011010001000",
				"011110011001",
				"011110011001",
				"010110000111",
				"011010001000",
				"100010101010",
				"011110011001",
				"100010001000",
				"100010011001",
				"011001100111",
				"011001111000",
				"011110011010",
				"011010011001",
				"011010101001",
				"011010111011",
				"011010101010",
				"011110101010",
				"011010011001",
				"011110101010",
				"100010101010",
				"100010011001",
				"010101000101",
				"010101010110",
				"011110011010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110011010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"100010111100",
				"100110111100",
				"100110101011",
				"100110011011",
				"100001111001",
				"011101101000",
				"011001101000",
				"011001101000",
				"010101100111",
				"010101010111",
				"011001010111",
				"011101101000",
				"011101100111",
				"100010001010",
				"011110001001",
				"011010001001",
				"011010101010",
				"010110011010",
				"010010101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010001000",
				"010110001001",
				"011010011001",
				"010110001001",
				"011010001001",
				"011110011010",
				"100010101011",
				"100010101011",
				"011110011010",
				"011010001001",
				"011010001000",
				"011010001000",
				"100010011010",
				"100110111011",
				"101010111011",
				"100110111011",
				"101010111011",
				"100110101011",
				"100010011001",
				"100010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110101010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"001101110111",
				"001110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010001110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001110111",
				"011001110111",
				"011001111000",
				"011001110111",
				"011001110111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001001000100",
				"001001000100",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001010101",
				"001101010101",
				"001101010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001000100",
				"001101000100",
				"001101000011",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001100110011",
				"001000110010",
				"000100100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"001100110011",
				"010101010101",
				"011001100110",
				"011101111000",
				"100010001001",
				"100110011001",
				"100110101010",
				"101010101011",
				"101010111011",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110101010",
				"100010101010",
				"100010111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010111100",
				"100010111011",
				"100010111011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010010001001",
				"010010001000",
				"010010001001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011001",
				"011010001000",
				"011010011000",
				"011010101001",
				"011110101001",
				"011110011001",
				"011010001000",
				"011110011001",
				"011110101010",
				"011010011000",
				"010110011000",
				"011110101010",
				"100010101010",
				"011110011000",
				"010101100111",
				"010101111001",
				"100010111101",
				"100010101100",
				"011010011010",
				"010010011000",
				"011011001010",
				"011010111010",
				"011010101010",
				"011010011001",
				"100110101010",
				"101010011010",
				"011001010110",
				"010001000101",
				"100010001001",
				"100010101011",
				"011110101011",
				"011010101011",
				"011010011010",
				"011110011010",
				"011110101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110101100",
				"011110101011",
				"011110101010",
				"100010011010",
				"011101111000",
				"100001111001",
				"100110001010",
				"101010011011",
				"101010101100",
				"101010101100",
				"100110101100",
				"100110101011",
				"100010011011",
				"100010011011",
				"100010011011",
				"011110001010",
				"011110011010",
				"011110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110011011",
				"011010011011",
				"011010011011",
				"011110011011",
				"011110011011",
				"011010011010",
				"011010011010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011000",
				"010010001000",
				"011110101010",
				"010101110111",
				"010101100111",
				"010101100111",
				"011110001001",
				"011110001001",
				"011110001001",
				"100010011010",
				"100110101011",
				"100010101011",
				"100010101011",
				"011110101010",
				"011110011001",
				"011110011001",
				"011110101010",
				"011110101010",
				"011110011001",
				"011010011010",
				"011010011001",
				"010110001001",
				"010010001000",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011000",
				"001110001000",
				"001110001000",
				"001110000111",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010101100110",
				"011001100111",
				"011001100110",
				"010001010101",
				"001100110100",
				"001000110011",
				"001000110011",
				"001000110100",
				"001101000100",
				"001101000101",
				"001101010101",
				"010001010101",
				"010001010101",
				"010001100110",
				"001101010101",
				"001101010100",
				"001001000100",
				"001001000100",
				"001101010101",
				"010001100110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101110110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010101100101",
				"010101100110",
				"010101100110",
				"010001010101",
				"001101000011",
				"000100100010",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"001100110100",
				"011001100110",
				"011101111000",
				"100010001000",
				"100010011001",
				"100110101010",
				"101010101011",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110101010",
				"100110101011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"010110101010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011001",
				"011010011001",
				"011010101001",
				"011110101001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011110101001",
				"011110101010",
				"011010101001",
				"011010011001",
				"011110101010",
				"100010101010",
				"011010001000",
				"010001110111",
				"010110001010",
				"100010111101",
				"100010101100",
				"011010011010",
				"010010011000",
				"010110111001",
				"010110111010",
				"011010101010",
				"100010101010",
				"100010011001",
				"011101100110",
				"010101000101",
				"011101100111",
				"100010011010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011010101010",
				"010110101011",
				"010010101011",
				"010110101100",
				"011010101011",
				"011010011011",
				"011010011010",
				"010101111000",
				"011110001000",
				"101010101010",
				"101110101100",
				"101110111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100010111100",
				"011110101100",
				"011110101011",
				"011110011011",
				"011110101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110011011",
				"010110011011",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101001",
				"010110011000",
				"011110101010",
				"011001110111",
				"010001000101",
				"011001111000",
				"100110101011",
				"100110111011",
				"100110111100",
				"100010101010",
				"011110011010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110001001",
				"011010101010",
				"011110101010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010101010",
				"010110011001",
				"010110101001",
				"010110101001",
				"010110011001",
				"010010011001",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011001111000",
				"001101000100",
				"000100010001",
				"000100010010",
				"001000100010",
				"000100010010",
				"001000110011",
				"001101000101",
				"010001010101",
				"010001100110",
				"010101100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110000111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"001101000100",
				"001000110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100100010",
				"001000010001",
				"001000010001",
				"001000010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100011",
				"010001000101",
				"011001100111",
				"011110001000",
				"100010011001",
				"100110011001",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010101010",
				"011110101010",
				"011010011001",
				"011010011001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110101010",
				"011110101001",
				"011010011000",
				"011010001000",
				"011110011001",
				"100010101010",
				"100010101010",
				"011110101010",
				"011010101001",
				"011110101010",
				"100010101010",
				"010101110111",
				"010001110111",
				"011010011010",
				"011110111100",
				"100010011100",
				"011110101011",
				"010010011000",
				"010110101001",
				"011110111010",
				"100010111011",
				"100110101011",
				"011101111000",
				"010001000101",
				"010101010110",
				"100010001001",
				"100010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111011",
				"010110101100",
				"011010101100",
				"011010011011",
				"011010001010",
				"011110011011",
				"011110001000",
				"011101110111",
				"101110101011",
				"101010111100",
				"100110111100",
				"100010111100",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010011011",
				"011010011011",
				"010110011011",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110101001",
				"011010101001",
				"011010101001",
				"100010111011",
				"100010011010",
				"010101010110",
				"011010001001",
				"011110011010",
				"011010011010",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110011000",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010101010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101001",
				"011010011001",
				"011010001000",
				"010101110111",
				"011001110111",
				"010101100110",
				"001101000100",
				"001101000100",
				"010101100110",
				"011110001000",
				"011110001000",
				"010101110111",
				"010110001000",
				"011010001001",
				"011010001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010110001000",
				"010110011000",
				"011010011001",
				"010110011000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010110000111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"011001110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001000100",
				"001000100010",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100010",
				"000100100010",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100010",
				"001101000100",
				"010101100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111011",
				"100110101011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110101010",
				"011110101010",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"100010111100",
				"100011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101100",
				"011010111100",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010101100",
				"010110101011",
				"010110011011",
				"010110101011",
				"010110101011",
				"011010101100",
				"011010111100",
				"011110111100",
				"011110111101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"011010011001",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010101001",
				"011010011000",
				"011010011001",
				"100010101010",
				"100010101010",
				"011110101001",
				"011110101001",
				"011110101010",
				"011110101010",
				"100010011001",
				"010101110111",
				"010001110111",
				"011010101011",
				"011110111100",
				"100010101011",
				"100010101011",
				"010110011001",
				"011010101001",
				"100010111010",
				"100110101011",
				"011101111000",
				"010101010110",
				"011001100111",
				"011110001001",
				"011110011001",
				"100010101011",
				"011010101011",
				"010110111100",
				"010110111011",
				"011010111011",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111011",
				"011010101011",
				"011010101100",
				"011110101100",
				"011110011011",
				"100110101011",
				"100010011001",
				"011101110111",
				"100110101010",
				"100010101011",
				"011110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"010010011010",
				"010010011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010010101010",
				"010010101010",
				"010010011001",
				"010110101001",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011001",
				"011110011001",
				"011001101000",
				"010101010111",
				"011110001001",
				"011010011010",
				"010110011001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"010010001001",
				"001101111000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010001111000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010001000",
				"011110011001",
				"100010101010",
				"011010001000",
				"001101000100",
				"010001010101",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010110001000",
				"010110011000",
				"010110011000",
				"010110011000",
				"010110011000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101010101",
				"001101000011",
				"000100100001",
				"000000000000",
				"000000010001",
				"000000010001",
				"000000010001",
				"000000010001",
				"000100010001",
				"000100100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100100001",
				"000100010001",
				"000000010001",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000000010001",
				"001000100010",
				"010001010101",
				"011001110111",
				"011110001000",
				"100010011001",
				"100110011001",
				"100110101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010101011",
				"100110101011",
				"100110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111011",
				"100010101011",
				"011110101010",
				"011110101010",
				"100010101011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110111100",
				"100010111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011110111101",
				"011010111101",
				"011010111101",
				"011110111101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"011010101100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010111011",
				"011010111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010111011",
				"011010101010",
				"011010011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110001001",
				"011110011010",
				"100010101011",
				"011110101010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110101010",
				"100010101010",
				"011110011001",
				"011010011000",
				"011010011001",
				"011110101010",
				"100010101010",
				"100010101010",
				"011001110111",
				"010110000111",
				"011010111011",
				"011110111011",
				"100010101011",
				"100010101011",
				"011010011001",
				"011110011001",
				"101010111011",
				"100010001000",
				"011001010110",
				"011001100111",
				"011110011010",
				"100010101011",
				"011110011010",
				"011110101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111010",
				"010110111010",
				"011010111010",
				"011010101010",
				"011110111011",
				"011010011010",
				"011110101011",
				"100010101100",
				"100110101011",
				"100010011010",
				"011001110111",
				"011110001000",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110011010",
				"011010011010",
				"011010101011",
				"011110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010101010",
				"011110111011",
				"011110101011",
				"100010101011",
				"100010011010",
				"011101111000",
				"011101100111",
				"011001010111",
				"011001000110",
				"011001000110",
				"100001111001",
				"100010001010",
				"011110011010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"011010001001",
				"011010001001",
				"010110001000",
				"010110001001",
				"010110011001",
				"010010001001",
				"010110101010",
				"010110101010",
				"010010011001",
				"010110101010",
				"011010111011",
				"011010101010",
				"010010011001",
				"001110001000",
				"010010001000",
				"010010001001",
				"010010011001",
				"010010001000",
				"001110001000",
				"010010011001",
				"010110011001",
				"010110001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001000",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001110111",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010101001",
				"010110011001",
				"010010001000",
				"010001110111",
				"001101110110",
				"001101110110",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010101110111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100101",
				"001101010101",
				"001101000100",
				"001101010100",
				"001101010101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001010101",
				"010001010100",
				"001101000100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001010100",
				"001101010100",
				"001101000100",
				"001101000011",
				"001000110010",
				"000100100010",
				"000100100001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100100010",
				"001100110100",
				"010101100110",
				"011001110111",
				"011110001000",
				"100010011001",
				"100110101010",
				"101010111010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100010101011",
				"100010101010",
				"100010101011",
				"100010111011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111011",
				"011110101011",
				"011110111011",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010101100",
				"011010101011",
				"011010101100",
				"011010111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"010110101011",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011111001101",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010111011",
				"010110101010",
				"010110011001",
				"010110011010",
				"011010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"100011001100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"011110101010",
				"100010111011",
				"011110101010",
				"010110011001",
				"011010011001",
				"011110101010",
				"100010101010",
				"011110101001",
				"011010011001",
				"011010011000",
				"011110011001",
				"100010111010",
				"100110111011",
				"100010101010",
				"010101110111",
				"010110001000",
				"011010111010",
				"011010111010",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110011001",
				"100110011001",
				"011001010110",
				"011001010110",
				"011110001010",
				"011110101011",
				"011110111100",
				"100010111100",
				"011110101011",
				"010110011010",
				"011010101011",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111010",
				"011010101010",
				"100010111100",
				"011010011010",
				"011110101010",
				"100010111011",
				"011110011010",
				"011010001001",
				"011010001000",
				"011010011001",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101100",
				"011010101011",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010101010",
				"011110011001",
				"011001100111",
				"010101000101",
				"010000100100",
				"010100100101",
				"011101000110",
				"011101000111",
				"100110001010",
				"101110111101",
				"100110011011",
				"011110011010",
				"011010101011",
				"010110011010",
				"010110101010",
				"010010011010",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110101010",
				"010110101010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011001",
				"011010101010",
				"010110011001",
				"010010011001",
				"010110011001",
				"011110011010",
				"011010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"000101000100",
				"000000100011",
				"000101000100",
				"010001110111",
				"011010011001",
				"011010011001",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011000",
				"010110011001",
				"010110011000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"001101010101",
				"001101010100",
				"001001000100",
				"001001000100",
				"001101010101",
				"010001010101",
				"010001100101",
				"010001100110",
				"001101010100",
				"001101010100",
				"001101010101",
				"001101010100",
				"001101010100",
				"001101010101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101100110",
				"010101110110",
				"011001110111",
				"011001110111",
				"011001110110",
				"010101100110",
				"010101010101",
				"010101100110",
				"010101110110",
				"011001110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010001100101",
				"001101000100",
				"001000110011",
				"001000110010",
				"000100100010",
				"000100100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000110011",
				"010001000100",
				"010101100110",
				"011101110111",
				"100010011001",
				"100110101010",
				"100110101010",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111100",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111100",
				"100010111100",
				"100010111101",
				"100011001101",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010101100",
				"011010101011",
				"011010111100",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"010110111100",
				"010110101011",
				"010110101100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110011010",
				"010010001001",
				"010110011010",
				"011010101011",
				"011110111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111011",
				"011010101010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011110101011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110101011",
				"011110101011",
				"011010011001",
				"010110011001",
				"011010101001",
				"011110101010",
				"011110101010",
				"011110011001",
				"011110011001",
				"011110011001",
				"011110101010",
				"100010111011",
				"100110111011",
				"011110011001",
				"010001100110",
				"011010001000",
				"011010111010",
				"011010101010",
				"011110101011",
				"100010101011",
				"100010111011",
				"011010001000",
				"011001010101",
				"011001000101",
				"011101111000",
				"100010011011",
				"011010101100",
				"011010111100",
				"100011001100",
				"011110111011",
				"010110001001",
				"011010011010",
				"011110101011",
				"011110111100",
				"011010111100",
				"011010111100",
				"011110111011",
				"011110101011",
				"011110101010",
				"100010111010",
				"100011001011",
				"011110101010",
				"010101100111",
				"010101100111",
				"011110011011",
				"100010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010101011",
				"011010011010",
				"011110101011",
				"100110111100",
				"101010111100",
				"100110101011",
				"100010001001",
				"011101111000",
				"011001100111",
				"010101010110",
				"010101010110",
				"010001000101",
				"010001000110",
				"010101000110",
				"011001101000",
				"100110001010",
				"100010001010",
				"100110011011",
				"101010111100",
				"100010101011",
				"011110101011",
				"011010111011",
				"010110101011",
				"010110111011",
				"010010101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"011010101010",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110101010",
				"011010101010",
				"010110001000",
				"010110001000",
				"011010001001",
				"011110101010",
				"011110101010",
				"011010011001",
				"011010001001",
				"010001110111",
				"010101110111",
				"010101111000",
				"010001110111",
				"001101100110",
				"001001010101",
				"001101110111",
				"011010011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"011010011001",
				"010010001000",
				"010110001000",
				"010110011001",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"010110001000",
				"010101110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010101110110",
				"010001100110",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101110110",
				"010001100110",
				"001101010101",
				"010001100101",
				"010001100110",
				"010101100110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101010101",
				"010001000100",
				"001000110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000100010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"001101000100",
				"010101010101",
				"011001110111",
				"100010001000",
				"100010011001",
				"100110101010",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101010111100",
				"101010111100",
				"101110111100",
				"101110111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110101011",
				"100010101011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100010111100",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100111001100",
				"100111001101",
				"101011001101",
				"101011001110",
				"100111001101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"011111001110",
				"100011001110",
				"011111001110",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010101100",
				"011010111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111001110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"010110111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110011010",
				"011010101011",
				"011110111100",
				"100011001101",
				"100011001100",
				"011110111100",
				"011110111011",
				"010110011010",
				"010010001001",
				"010110011001",
				"011010101010",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101010",
				"010110011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110101001",
				"011110101010",
				"100010111011",
				"100010101010",
				"100010111011",
				"100010101010",
				"011010001000",
				"010001010101",
				"011010011001",
				"011110111010",
				"010110101001",
				"011010101010",
				"011110101011",
				"100010111011",
				"010101100110",
				"001100010010",
				"011101010110",
				"100010011010",
				"011110101011",
				"011010101100",
				"011010111101",
				"011110111100",
				"011110111011",
				"011010101010",
				"011010101010",
				"011110101011",
				"011110111100",
				"011110111101",
				"011010111100",
				"011110101100",
				"100010111011",
				"100010101010",
				"100111001011",
				"011110101000",
				"010001110110",
				"010101100110",
				"100010011010",
				"100110111101",
				"011110101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011010011010",
				"011110011010",
				"100010011010",
				"100010001001",
				"011101101000",
				"011001010110",
				"011001000110",
				"011001010110",
				"011101100111",
				"011101111000",
				"011110001000",
				"011110011010",
				"100010011010",
				"100010101011",
				"100110111100",
				"100010011011",
				"100110111100",
				"100010101011",
				"011110101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"010110111011",
				"010110101011",
				"010010101010",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010011010",
				"011110101011",
				"011110101011",
				"010110101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010010011001",
				"010010001000",
				"011010011001",
				"011010001001",
				"010001100111",
				"010001010110",
				"010101100110",
				"010001010110",
				"001101000101",
				"010101111000",
				"010001100110",
				"001101100110",
				"010001111000",
				"010110001000",
				"010010001000",
				"010110001000",
				"011010011001",
				"010110001001",
				"011010011010",
				"010110001001",
				"010110001000",
				"011010011010",
				"010110011001",
				"010010001001",
				"010110011001",
				"010001111000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010001110111",
				"010101110111",
				"011010001000",
				"010110001000",
				"010101110111",
				"010001100111",
				"001101100110",
				"001001010101",
				"001101010101",
				"001101100101",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010101110111",
				"010101110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101110111",
				"011001110111",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001000100",
				"001000110010",
				"000000010001",
				"000000010001",
				"000100100010",
				"001000110011",
				"001100110011",
				"001000110011",
				"001000100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100100001",
				"000100100010",
				"000100010001",
				"000000010001",
				"000000010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"001000100010",
				"010001000100",
				"010101100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"011110101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011110111100",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"011010101011",
				"010110011010",
				"010010001001",
				"010110011010",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101010",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"011110101010",
				"011110101011",
				"100010111011",
				"011110101010",
				"011010011001",
				"011110101010",
				"100010101010",
				"100010101010",
				"100110111011",
				"011110011001",
				"010001100110",
				"010001100110",
				"011010011001",
				"011110111010",
				"011010111010",
				"011010111011",
				"010110101010",
				"011110101010",
				"011110011001",
				"010000110011",
				"011001010110",
				"100010101011",
				"011110111100",
				"011010101101",
				"011010111101",
				"011010101011",
				"011110111011",
				"011111001011",
				"010110101010",
				"010110001001",
				"011110111100",
				"100011001101",
				"011110111100",
				"100010111100",
				"100110111100",
				"100110111011",
				"011110011000",
				"010001100101",
				"010001100101",
				"011001111000",
				"100110011011",
				"100110101100",
				"100010101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"011110111100",
				"011110101010",
				"010101110111",
				"010101100111",
				"011001010111",
				"011101010110",
				"100101101000",
				"101010001010",
				"100110001001",
				"100110101010",
				"100010101010",
				"011110101010",
				"011010111011",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111011",
				"010010101010",
				"010010011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010010001001",
				"011010001010",
				"011010011010",
				"011010011010",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010011001",
				"011010001001",
				"010101110111",
				"001101000101",
				"010001000101",
				"100001111000",
				"011101111000",
				"011110011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"011010011001",
				"011010101010",
				"011010011010",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010001111000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110110",
				"010001100110",
				"010001100110",
				"010101110110",
				"011001110111",
				"011001110111",
				"011001110111",
				"010101110110",
				"010001100101",
				"010001100101",
				"010101100110",
				"010101100110",
				"010001100101",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001010101",
				"001101010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101010101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101100110",
				"010101100110",
				"010001010101",
				"010001000100",
				"001101000100",
				"001000110011",
				"000100100010",
				"000100100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"001000110011",
				"010001010101",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101010111011",
				"101010111011",
				"100110111011",
				"100110111011",
				"100110111100",
				"101010111100",
				"101010111100",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111101",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"010110011010",
				"011010101011",
				"011110111100",
				"100011001100",
				"011110111100",
				"011110111011",
				"011010101010",
				"010110011010",
				"011010101010",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110111011",
				"100010111011",
				"011110101010",
				"011110101010",
				"100010111011",
				"100010101010",
				"100010101010",
				"100010101011",
				"011110011001",
				"010001100111",
				"010101111000",
				"100010101010",
				"011110101001",
				"011010101001",
				"011111001011",
				"011010111011",
				"100010111011",
				"011010001000",
				"010000110011",
				"011001100111",
				"011110111011",
				"011010111100",
				"011010111101",
				"011010111101",
				"011010101011",
				"011010111011",
				"011111001100",
				"011010101010",
				"011010011010",
				"011110101011",
				"011110111100",
				"100010111100",
				"100110111100",
				"011110011010",
				"010101110111",
				"010101110111",
				"011010001000",
				"011110011001",
				"100110101011",
				"100110011011",
				"100010011011",
				"100010101100",
				"011110111101",
				"011110111100",
				"011010101100",
				"011010101100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011110101011",
				"011010001001",
				"010101100111",
				"011001100111",
				"100101111001",
				"101010001010",
				"101010001010",
				"100110011010",
				"100010101010",
				"011110101010",
				"010110111010",
				"010010111010",
				"010010111011",
				"010010111011",
				"010010111011",
				"010010101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010011011",
				"011010011010",
				"011010101011",
				"010010011010",
				"010010101010",
				"010110101011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010110011010",
				"011010011011",
				"011010011011",
				"011010011010",
				"011010011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101001",
				"010110011001",
				"011110101010",
				"100010101010",
				"100010011010",
				"011001100111",
				"011001010111",
				"100001111001",
				"100010001010",
				"011010001001",
				"011010011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110001001",
				"010001111000",
				"010001111000",
				"010010001001",
				"011010011010",
				"010010001000",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010101110111",
				"010110000111",
				"010101110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010101110110",
				"010101110111",
				"010101110110",
				"001101010100",
				"001001000100",
				"001001000100",
				"001001000011",
				"001001000011",
				"001001000100",
				"001101000100",
				"001101010100",
				"001101010100",
				"001101010101",
				"010001100101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010101100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"011001110111",
				"010101010101",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001000100010",
				"000100100010",
				"000100100001",
				"000100010001",
				"000000010001",
				"000000010000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"100111001101",
				"100110111100",
				"100110111100",
				"100010111100",
				"100010111100",
				"100011001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"010110011010",
				"011010101010",
				"011110111011",
				"100011001101",
				"100011001101",
				"011111001100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011010101010",
				"011110101010",
				"100010111011",
				"100010111011",
				"100010101011",
				"100010101010",
				"011110011001",
				"011010011001",
				"100010101011",
				"100010111011",
				"011110101010",
				"011110111011",
				"011111001100",
				"011010111010",
				"100111001100",
				"011010001000",
				"001100110011",
				"011001111000",
				"011010111011",
				"010110111100",
				"011010111101",
				"011110111101",
				"011010101011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011010011010",
				"100010101011",
				"101011011101",
				"100010111011",
				"011001111000",
				"010101100111",
				"010101110111",
				"011010001001",
				"011110101011",
				"100010111100",
				"100110111100",
				"101010111101",
				"100010101100",
				"011110011011",
				"011110101100",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"011010111010",
				"010110001000",
				"010101100111",
				"100010011010",
				"100110101011",
				"100010011010",
				"100110111011",
				"011110101011",
				"011010111011",
				"010110111011",
				"010010111011",
				"010110111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"100010101100",
				"011110011011",
				"011010011010",
				"011010011011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"011010101011",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"100010101011",
				"100010101010",
				"011110001001",
				"011110001000",
				"011001111000",
				"011001100111",
				"011001111000",
				"011001111000",
				"011010011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"010110011010",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010010001000",
				"001110001000",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101111000",
				"010001100110",
				"010101110111",
				"010101110111",
				"010001100111",
				"010001110111",
				"010110001000",
				"010110001001",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110000111",
				"010110000111",
				"010001110111",
				"010001100110",
				"010001110110",
				"010101110111",
				"010001110110",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110111",
				"010001100110",
				"001101010101",
				"000100110011",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001010101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000100",
				"001101000011",
				"001100110011",
				"001000110010",
				"001000100010",
				"000100100001",
				"000100010001",
				"000100010001",
				"000100010001",
				"000100010000",
				"000100000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"100111001100",
				"100111001100",
				"101010111100",
				"101010111100",
				"100110111100",
				"100110111011",
				"100010111011",
				"100010111011",
				"100010111100",
				"100111001100",
				"100111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001100",
				"100111001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100110111101",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111001110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101100",
				"010110011011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110111011",
				"100011001100",
				"100111001101",
				"100011001100",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"011110101011",
				"011010101010",
				"011110101010",
				"100010111011",
				"100010101011",
				"100010101010",
				"100010101010",
				"011110101010",
				"100110111100",
				"100111001100",
				"011110101011",
				"100010111011",
				"100011001100",
				"011010111011",
				"011010111010",
				"100111001011",
				"010101100110",
				"001101000100",
				"011110001001",
				"011010111100",
				"010110111100",
				"011110111101",
				"011110111101",
				"011010101011",
				"011010111011",
				"011010111100",
				"100010111100",
				"011010011010",
				"011010001001",
				"100010011010",
				"011001110111",
				"010101100110",
				"011001111000",
				"100010101011",
				"100010111100",
				"100010111101",
				"011110101100",
				"100010111100",
				"100111001101",
				"100111001101",
				"011110101011",
				"010110101010",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010111010",
				"011110111011",
				"010110001000",
				"010001100111",
				"011110011001",
				"100010101011",
				"011110101011",
				"011110111100",
				"011010101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110101011",
				"100010101100",
				"011110101011",
				"011010011011",
				"010110011010",
				"010110101011",
				"011010101011",
				"010110101011",
				"011010101010",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110011010",
				"010110101011",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110011010",
				"100010011010",
				"100010101010",
				"100010001001",
				"011001100111",
				"010001000101",
				"010001000101",
				"011001110111",
				"011001111000",
				"011010001001",
				"011010001001",
				"011010011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110101010",
				"011010101011",
				"011010101010",
				"010110011001",
				"001110001000",
				"010010011001",
				"010010001000",
				"010010011001",
				"010110011001",
				"010010011001",
				"010010001000",
				"010010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010001100110",
				"010101110111",
				"010101110111",
				"010001110111",
				"010101111000",
				"010110001001",
				"010110001001",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"011010011000",
				"010110000111",
				"010001100110",
				"010001110110",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010101110110",
				"010001110110",
				"010001100110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"001101010101",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101010101",
				"010001010101",
				"010001010101",
				"010101010101",
				"010001000100",
				"010001000011",
				"001100110011",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000110010",
				"001000110010",
				"001100110011",
				"001100110011",
				"001100110011",
				"001100110010",
				"001000100010",
				"000100010001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001110",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011110111100",
				"011111001101",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011110111011",
				"011110111100",
				"100011001100",
				"100011001101",
				"100011001101",
				"011110111100",
				"010110101010",
				"011010101010",
				"011110111011",
				"100011001100",
				"100010111100",
				"100010111011",
				"011110101010",
				"011110111011",
				"100010111100",
				"011110101011",
				"011110011010",
				"011110011010",
				"011110101011",
				"100111001101",
				"100111001101",
				"011110111100",
				"100010111100",
				"011110101011",
				"011110111011",
				"100111001100",
				"100010101001",
				"001101000011",
				"010001010101",
				"011110011010",
				"011011001100",
				"010110111100",
				"011110111101",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"100010101011",
				"011110001000",
				"001101000100",
				"010101010101",
				"100110011010",
				"100010011011",
				"100010111100",
				"011110111101",
				"011110111101",
				"011111001110",
				"011010111101",
				"011010111011",
				"011110111100",
				"100011011101",
				"011010111011",
				"010110101011",
				"011010111100",
				"011111001100",
				"010110111100",
				"011010111100",
				"011011001101",
				"010110111100",
				"010111001100",
				"010110111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110101010",
				"011010111011",
				"100010111011",
				"100110111011",
				"011110011001",
				"010101100111",
				"010101111000",
				"011110101011",
				"100010111100",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101011",
				"010110101011",
				"010010101010",
				"010010101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010010011010",
				"010110101010",
				"011010111100",
				"011010111011",
				"011010101010",
				"011010101010",
				"011110101011",
				"100010111100",
				"011110101100",
				"011110101011",
				"100010101011",
				"100110111100",
				"100110101011",
				"100001111001",
				"011001010110",
				"011101010111",
				"011001010110",
				"010101000101",
				"011001010110",
				"011110001001",
				"011110011001",
				"011110011010",
				"011110101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"001110001000",
				"001101110111",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"011010001001",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101111000",
				"011010001001",
				"011010001000",
				"011010001000",
				"011010001001",
				"011010011001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010101110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"011010000111",
				"011001110111",
				"010101100110",
				"001101010101",
				"001101010100",
				"001001000100",
				"000100110011",
				"001101000100",
				"001101000100",
				"001101010100",
				"001101010101",
				"010001100101",
				"010001100110",
				"010101100110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010001000100",
				"001101000011",
				"001100110011",
				"001000110010",
				"001000100010",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010101",
				"010101010100",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001010100",
				"010001010100",
				"010001010100",
				"001101000100",
				"001100110011",
				"001000100010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010001001",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010111011",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111100",
				"100111001100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100110111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"100111011101",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011001110",
				"101011001110",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111001101",
				"100111001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100011011101",
				"100011011101",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011111001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011110111100",
				"011010101100",
				"011010101100",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111100",
				"100011001101",
				"100011001101",
				"100010111101",
				"011110111100",
				"011110111100",
				"011110101011",
				"011110111100",
				"011110111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100011001100",
				"100011001100",
				"011110111011",
				"010110101011",
				"011010111011",
				"100011001100",
				"100111001101",
				"100111001100",
				"100010111100",
				"011110111011",
				"011110111011",
				"100010111100",
				"011110101010",
				"011010001001",
				"011110011010",
				"100010101011",
				"100111001101",
				"100011001100",
				"011110111100",
				"011110111101",
				"011110111100",
				"101011011101",
				"100110111010",
				"010101010101",
				"001101000011",
				"011001110111",
				"100010101011",
				"011011001100",
				"010110111100",
				"011010111100",
				"011110101100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101010",
				"100010111011",
				"100010011001",
				"010101000101",
				"011001010110",
				"101010101011",
				"100110101011",
				"011110101100",
				"011110111101",
				"011010111110",
				"011011001110",
				"010110111100",
				"010110111011",
				"011010111011",
				"011111001100",
				"011111011101",
				"010010101010",
				"010110101010",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"010110111100",
				"011011001101",
				"011011001101",
				"010110111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"100010111011",
				"100010001001",
				"010101010110",
				"010101100110",
				"100010011010",
				"100010111100",
				"011110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010101100",
				"011010101011",
				"011110101011",
				"011110101011",
				"011010101010",
				"010110101010",
				"010010101010",
				"010010011010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111100",
				"010110101010",
				"010110101010",
				"011110111100",
				"100011001101",
				"100011001100",
				"100010111100",
				"100010111100",
				"100010101100",
				"100010111100",
				"100010101011",
				"100010011010",
				"011110001010",
				"100010011010",
				"101010011011",
				"101110101011",
				"101010011010",
				"101010011010",
				"100110001001",
				"100110011010",
				"100110101011",
				"011110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001000",
				"010010011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010011001",
				"010010001000",
				"010001111000",
				"010001111000",
				"001101100111",
				"001101100110",
				"001101010110",
				"001101100110",
				"010001110111",
				"010101110111",
				"011110011001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010011010",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"010101110111",
				"001101010101",
				"001001000100",
				"001001000101",
				"001001000100",
				"001001000100",
				"001001000100",
				"001001010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010110000111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110111",
				"010101110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"001101000100",
				"001001000011",
				"001001000100",
				"001101010101",
				"010001010101",
				"001101010100",
				"010001100110",
				"010101110110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010001010100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101100101",
				"010001010101",
				"010001010100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"001000100011",
				"001101000100",
				"010101010101",
				"011001100111",
				"011101111000",
				"100010001001",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111100",
				"100110111011",
				"100110111011",
				"100110111100",
				"100111001100",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011001110",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111011110",
				"100111001110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011111001101",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011110111101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111011",
				"010110101011",
				"011010101011",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011110111100",
				"100011001100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100010111100",
				"011110111100",
				"011110111011",
				"011110111100",
				"011111001100",
				"100011011101",
				"100111001101",
				"100110111100",
				"100010111011",
				"011110111011",
				"011110111011",
				"100011001100",
				"011110011010",
				"011010001001",
				"100010101011",
				"100110111100",
				"100011001101",
				"011110111011",
				"011010101011",
				"011010111100",
				"100010111101",
				"101011001100",
				"011110001000",
				"010101010100",
				"010101010101",
				"011110001001",
				"100010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111011",
				"011111001100",
				"011010111011",
				"011110111010",
				"011110101010",
				"011001100111",
				"011001010111",
				"100010011010",
				"100110111100",
				"011110111100",
				"011111001101",
				"011010111101",
				"010110111100",
				"010110111100",
				"011011001101",
				"011110111100",
				"011010101011",
				"011111001100",
				"011010111011",
				"010110101010",
				"011010101011",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010101011",
				"100010111100",
				"100110111100",
				"100010011010",
				"011001110111",
				"011001010110",
				"010101000101",
				"011001111000",
				"100010101011",
				"011110101011",
				"011010101011",
				"011010111100",
				"011111001101",
				"011010111101",
				"011110111100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111011",
				"011010101011",
				"011110101011",
				"011110101011",
				"100110111100",
				"100110111100",
				"100010101011",
				"011110011010",
				"011110001010",
				"011010001001",
				"011110011010",
				"100110111100",
				"101111011101",
				"101111011101",
				"101011001100",
				"101011001100",
				"101010111100",
				"100110101010",
				"100110101011",
				"100110111011",
				"100010101010",
				"011110011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"011010001001",
				"010001100111",
				"001001000100",
				"001001000100",
				"001001000101",
				"001101010101",
				"001101100110",
				"001101100110",
				"001101100111",
				"010001111000",
				"011010001001",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001001",
				"011010011001",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"001101010101",
				"000100110011",
				"000100110011",
				"001001000100",
				"001101100110",
				"010001110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"001101110111",
				"010001110111",
				"010010001000",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010101110110",
				"010001100110",
				"001101010101",
				"001101010100",
				"001101010101",
				"010001100101",
				"010001100101",
				"001101100101",
				"001101010101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010101110110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000011",
				"001101000100",
				"010001010100",
				"010101100101",
				"010101100101",
				"010101100101",
				"010101010101",
				"010101010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010101",
				"010001010101",
				"010001010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000110011",
				"010001000101",
				"010101010110",
				"011001110111",
				"011110001000",
				"100010001000",
				"100110011001",
				"100110101001",
				"101010101010",
				"101010111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"101111001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101011001100",
				"101011001100",
				"101010111100",
				"101010111011",
				"100110111011",
				"100110111011",
				"101011001100",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"101011001110",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111011101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"011111011111",
				"011111011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011001110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"100011001101",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011010111100",
				"011010101011",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101011",
				"011010101011",
				"011110101011",
				"100011001100",
				"100011001101",
				"100011001100",
				"100011001101",
				"100011001101",
				"011110111011",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011011101",
				"100111011101",
				"100111001100",
				"100010101011",
				"011110101010",
				"011110111011",
				"011110111100",
				"100011001100",
				"011110101010",
				"011010001001",
				"100010101011",
				"100111001100",
				"011110111100",
				"011110111100",
				"011010111011",
				"100011001101",
				"100111001110",
				"100110111100",
				"100110101010",
				"101010101010",
				"011101110111",
				"100010011010",
				"100010101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011111001100",
				"011011001100",
				"010111001011",
				"011010111011",
				"100011001100",
				"100110111011",
				"011001010110",
				"011001100111",
				"100010101011",
				"011110101011",
				"011110111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011110111100",
				"011110101011",
				"011010101011",
				"100011001101",
				"011110111100",
				"010110011010",
				"011010111100",
				"011111001101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011110111101",
				"100111001101",
				"100111001101",
				"100010101011",
				"011001111000",
				"010101100111",
				"010101010110",
				"011001010110",
				"011101100111",
				"100010001001",
				"100010101010",
				"011010011010",
				"011010101011",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010101100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010010011010",
				"010110101010",
				"011010101011",
				"011110101011",
				"011110011010",
				"010101111000",
				"010101100111",
				"011001111001",
				"011110001010",
				"100010011011",
				"100110101100",
				"101010111101",
				"100110111100",
				"100010111100",
				"100010111011",
				"100010111011",
				"011110101010",
				"011010011010",
				"011110101010",
				"011010011001",
				"011110101010",
				"011110101010",
				"011010011010",
				"011110101010",
				"011010011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010010011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011010",
				"010010011001",
				"010110011010",
				"011010011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011010001001",
				"010001100110",
				"001000110100",
				"001101000100",
				"010101100111",
				"011010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010101111000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010110001000",
				"011010011000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010001110111",
				"010010000111",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010001100101",
				"001101000100",
				"001000110011",
				"001000110011",
				"001000110011",
				"001101000100",
				"001101000100",
				"010001010101",
				"010001010101",
				"010101100101",
				"010101100110",
				"010101110110",
				"010001100101",
				"010101100101",
				"010101100110",
				"010101100110",
				"010101100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"010001010100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"010001000100",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101010111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"100111001101",
				"101011011101",
				"101011011101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011101",
				"100111001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011110111101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111001110",
				"011110111101",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011101",
				"011111011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011010101011",
				"010110011010",
				"011010011011",
				"100010111100",
				"100011001101",
				"100011011101",
				"100011001101",
				"011111001100",
				"011110111011",
				"011110101011",
				"100011001101",
				"011110111100",
				"100011001101",
				"100111011110",
				"101011001101",
				"100010101011",
				"100010011010",
				"100010101011",
				"100010111011",
				"100011011101",
				"011111001100",
				"011010101010",
				"011110101010",
				"100010111100",
				"011111001100",
				"011110111100",
				"100010111100",
				"011010011011",
				"100110111101",
				"100111001101",
				"100010111100",
				"100111001100",
				"110011101110",
				"100110111100",
				"100010011011",
				"011110011011",
				"011110111101",
				"011010101100",
				"011110111100",
				"011010111100",
				"010110111100",
				"010111001011",
				"010111001011",
				"011010111011",
				"100111001100",
				"100110111011",
				"011001100111",
				"011001111000",
				"010110011001",
				"011011001100",
				"010111001100",
				"011010111101",
				"011110111101",
				"100010111101",
				"011110111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"100010111100",
				"011110111011",
				"011110111100",
				"011010111011",
				"011010101011",
				"011110111011",
				"100111011110",
				"100111001101",
				"100011001101",
				"100010111100",
				"100010101011",
				"011110001001",
				"010101010111",
				"010101000110",
				"011101101000",
				"100110001010",
				"101110101100",
				"100110011011",
				"100010011010",
				"011110101010",
				"011010101010",
				"010110101010",
				"011010101011",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010101100",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111011",
				"010110101011",
				"011010101010",
				"011010011010",
				"011110011010",
				"100110011011",
				"011101111001",
				"010001010110",
				"100010011011",
				"100110111100",
				"100110111100",
				"100010101100",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010101010",
				"010110101010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101011",
				"011110111011",
				"011010101011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010010011010",
				"010110101011",
				"010110101010",
				"010010011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110001000",
				"011010001000",
				"100110101011",
				"100010011010",
				"011001100111",
				"011001100111",
				"011001100111",
				"011110001000",
				"010110001001",
				"010010011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010110011000",
				"010110011000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110000111",
				"010110001000",
				"010110000111",
				"010001110111",
				"011110011001",
				"010101110111",
				"001101100101",
				"001101100110",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010001000",
				"001110000111",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"001110000111",
				"001110000111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001111000",
				"011001111000",
				"011001110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100110",
				"010101110111",
				"010101110110",
				"010101110110",
				"010101110110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010101100101",
				"010101100110",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001010101",
				"010001100101",
				"010001100101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001100101",
				"010101100110",
				"010001100101",
				"001101010100",
				"001101000100",
				"001101010100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001100110011",
				"010001000100",
				"011001100110",
				"011001110111",
				"011101111000",
				"100010001001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001011",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101010111100",
				"100110111100",
				"100110111100",
				"100111001100",
				"101011001101",
				"101011011101",
				"101011011110",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011001101",
				"100111001101",
				"100111001110",
				"100111001110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111001101",
				"011010111100",
				"011010101100",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100010111101",
				"011110111101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111001100",
				"011010101011",
				"011010011011",
				"011110101011",
				"100010111100",
				"100011001101",
				"100011011101",
				"011111001101",
				"011110111100",
				"011110111011",
				"100010111100",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111001101",
				"100111001101",
				"100110111100",
				"100110101011",
				"100010101011",
				"100011001100",
				"100011011101",
				"011111001100",
				"011010111011",
				"011110111011",
				"100010111100",
				"011111001100",
				"011111001100",
				"100010111100",
				"011110011010",
				"100110111101",
				"100010111100",
				"011110111100",
				"100011001101",
				"101011011110",
				"101011001110",
				"011010001010",
				"011110001011",
				"100010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"010111001011",
				"011111001011",
				"101011001100",
				"100010001001",
				"010001000101",
				"011010001001",
				"011111001100",
				"010111001100",
				"011011001101",
				"011010111101",
				"011110111101",
				"011110101100",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011110111011",
				"011110101010",
				"100110111100",
				"100110101011",
				"011110001001",
				"011010001001",
				"010101100111",
				"010001010111",
				"011001010111",
				"100001111001",
				"100110011011",
				"100110101011",
				"100110101100",
				"100110111101",
				"100111001101",
				"100111001100",
				"011110111011",
				"010110101010",
				"011010101010",
				"011110111100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"010110111011",
				"011010111011",
				"011010101010",
				"011110011010",
				"100010011010",
				"100010011010",
				"011001111001",
				"100110011011",
				"101010111101",
				"100010101100",
				"011110101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011110111011",
				"011010101011",
				"010110011010",
				"010010011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110011010",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011110101010",
				"011110011001",
				"011001111000",
				"010001010101",
				"010001000101",
				"010101010110",
				"011001100111",
				"010101110111",
				"010110001001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110011000",
				"010110011000",
				"010110011000",
				"010110011000",
				"010110001000",
				"010110000111",
				"010110001000",
				"011010001000",
				"011010011000",
				"011010011000",
				"011010011000",
				"010110001000",
				"010101110111",
				"001101010101",
				"001001000100",
				"001001000100",
				"001101010110",
				"010001110111",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"001110000111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011110001001",
				"011110001000",
				"011010001000",
				"010101100110",
				"001101010101",
				"001001000100",
				"001001000100",
				"001101010100",
				"001101010101",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110111",
				"010101110110",
				"010001100101",
				"001101000100",
				"010001010101",
				"010001010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010001010101",
				"001101000100",
				"001101010100",
				"010001010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101110111011",
				"101010111011",
				"101010111011",
				"101010111100",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101010111100",
				"100110111100",
				"100111001100",
				"101011001101",
				"101011011101",
				"101011011110",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101011011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011111",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001110",
				"100011001101",
				"100011001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111001110",
				"011110111101",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111001101",
				"011010111100",
				"011010101011",
				"011010101011",
				"011110111100",
				"100011001101",
				"100011011110",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011110111100",
				"011110111100",
				"100010111101",
				"100011001101",
				"100011001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011110111100",
				"011110101100",
				"100010111100",
				"100011001101",
				"100011011101",
				"011111001101",
				"011111001100",
				"011010101011",
				"011110101011",
				"100010111100",
				"100011001101",
				"100111011110",
				"100111011110",
				"100011001100",
				"100010111100",
				"100110111100",
				"100110111100",
				"100110111100",
				"101011011101",
				"100011001100",
				"011110111011",
				"011010101010",
				"011110111011",
				"011110111100",
				"011111001100",
				"011111001100",
				"100010111101",
				"011110011010",
				"100010101011",
				"011110101011",
				"011110111100",
				"011111001101",
				"100011001101",
				"101011011110",
				"011110001011",
				"010101111001",
				"011010101011",
				"011110111100",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011110111011",
				"100111001100",
				"100110011010",
				"011101101000",
				"011001101000",
				"100010101011",
				"011110111100",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111100",
				"011010111100",
				"011011001100",
				"011111001100",
				"011010101010",
				"010001010110",
				"011001010110",
				"011101100111",
				"010101000110",
				"011001100111",
				"011001111001",
				"011010001001",
				"011110011011",
				"100010111100",
				"100010111101",
				"011110111100",
				"011110101100",
				"100010111100",
				"100010111100",
				"100011001100",
				"100010111100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"011010111011",
				"010110101011",
				"011010111011",
				"011110101100",
				"011110101011",
				"011110011011",
				"011110101011",
				"011110111011",
				"011011001100",
				"010110111010",
				"011010111011",
				"011010111010",
				"011110101011",
				"100110111100",
				"100010001010",
				"011101101001",
				"100010001010",
				"011110011011",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101010",
				"011010011010",
				"011110101011",
				"011110111100",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010011010",
				"011110101011",
				"011110101010",
				"011010011001",
				"011010011010",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011110011010",
				"011110011001",
				"010001100111",
				"001101010101",
				"000100100011",
				"001000110100",
				"010101100110",
				"010101100111",
				"010101110111",
				"011010001001",
				"010110001001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"001101110111",
				"010001110111",
				"010110001000",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010001001",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100111",
				"010101111000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101100111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001010101",
				"010001010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110110",
				"010101110110",
				"010101110110",
				"010101100110",
				"010101110110",
				"010101100110",
				"010001100110",
				"010101100110",
				"010101100110",
				"010101100110",
				"010001100101",
				"010001010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111100",
				"101110111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101010111100",
				"101010111100",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011101",
				"101011011101",
				"101011011110",
				"100111011110",
				"100111011101",
				"100111001101",
				"101011001101",
				"100111001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001101",
				"011110111101",
				"011111001101",
				"100011001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010101011",
				"011010101011",
				"011110111100",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011010111011",
				"011010101011",
				"011110111100",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100010111101",
				"100111001101",
				"100111001101",
				"100011011101",
				"100011011101",
				"011111001100",
				"011010101011",
				"011110111011",
				"100011001101",
				"100011001101",
				"100111011110",
				"100011001101",
				"011110111100",
				"011110111100",
				"100111001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"100010111011",
				"011010011010",
				"011010011010",
				"011110111011",
				"011110111100",
				"011011001100",
				"011111001100",
				"100111001101",
				"011110011010",
				"011001111001",
				"010110011010",
				"011111001100",
				"011111011101",
				"011110111100",
				"100111001101",
				"100110101100",
				"010101101000",
				"010110001001",
				"011111001101",
				"011111001101",
				"011011001100",
				"100011001101",
				"100010111100",
				"100111001100",
				"100110101010",
				"100001111000",
				"100010001010",
				"101010101100",
				"101011001110",
				"011110101100",
				"100010111101",
				"011110111100",
				"011110111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011111001101",
				"010110101100",
				"010010101011",
				"011010111100",
				"100010111100",
				"011001110111",
				"010000110100",
				"011001000101",
				"011101100111",
				"100010011010",
				"100010111011",
				"011110111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011110111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011110111100",
				"011111001100",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010111001100",
				"010110111011",
				"011010111100",
				"011010101011",
				"011010011011",
				"011110011011",
				"100010101011",
				"100010101100",
				"011110111011",
				"011010111011",
				"010110111010",
				"011010111011",
				"011111001011",
				"011110101010",
				"100010101011",
				"011110001001",
				"011001101000",
				"011110001010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010101010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"011010101010",
				"010110011010",
				"011010101010",
				"011110101011",
				"011110101010",
				"011010011010",
				"011010011010",
				"011110101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110001000",
				"010001100111",
				"001101010110",
				"001101010101",
				"001101000101",
				"001000110100",
				"010001100111",
				"011010001001",
				"010101111000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011010011001",
				"010101111000",
				"010001100111",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010101100111",
				"011001111000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101110111",
				"010001110111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010110000111",
				"010001110111",
				"010010000111",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010101100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"001101100101",
				"001101010101",
				"010001100101",
				"010001100110",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010101100110",
				"010101110110",
				"010101100110",
				"010001010101",
				"001101010100",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101100110",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"100111001101",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101111011111",
				"101111101111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011001101",
				"100111001101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011111001101",
				"100011011110",
				"100011001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011101",
				"100011001101",
				"011110111100",
				"011010101011",
				"011010101011",
				"011110111100",
				"100011001101",
				"100111011101",
				"100111011110",
				"100011011110",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111001110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011110111100",
				"011111001101",
				"100111011110",
				"100111001110",
				"100111001110",
				"100011001101",
				"011111001100",
				"100011001101",
				"100111001101",
				"100111001101",
				"101011001101",
				"100111001100",
				"011110101010",
				"010110001001",
				"011010011010",
				"100010111100",
				"100011001101",
				"011011001100",
				"011111001100",
				"100111001101",
				"011110011011",
				"010001101000",
				"010110011010",
				"011111011101",
				"011011011101",
				"011111001100",
				"100011001101",
				"101010111101",
				"010101111001",
				"010010001001",
				"011111001100",
				"011111001101",
				"011010111100",
				"100011001101",
				"101011001101",
				"101010111100",
				"011110001001",
				"100110001010",
				"110010111110",
				"101010111110",
				"100110111110",
				"100110111110",
				"100010101101",
				"011110111100",
				"011110111100",
				"011011001100",
				"010111001100",
				"011011011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"011110111101",
				"011111001101",
				"011111001100",
				"100111001100",
				"100010101010",
				"010001000100",
				"011001010110",
				"100110101010",
				"100010101011",
				"011010111011",
				"010110111100",
				"010110111100",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"010111001100",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110111011",
				"011110111011",
				"100111001100",
				"100010101011",
				"100110101010",
				"011110001001",
				"011001100111",
				"011101111001",
				"011110001001",
				"100010101011",
				"011110101100",
				"011110101100",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010010101010",
				"010010101010",
				"011010111010",
				"011010111010",
				"011010101010",
				"010110011001",
				"010110011001",
				"011010101010",
				"011110111011",
				"100010111100",
				"011110101011",
				"011010011010",
				"010110001001",
				"001101100111",
				"001101100111",
				"010001100111",
				"010101111000",
				"011010001001",
				"011110001001",
				"011110011001",
				"011110011001",
				"011110011010",
				"011010011001",
				"010110011001",
				"011010011010",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"011010011001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101100111",
				"001101010110",
				"001101010101",
				"001001010110",
				"001101100110",
				"001101110110",
				"010001110111",
				"010010000111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110000111",
				"010110000111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110110",
				"010101110111",
				"010101110111",
				"011010001000",
				"011001110111",
				"010101110111",
				"010101100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101100101",
				"010001100110",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100101",
				"010001100110",
				"010001100110",
				"010101100110",
				"010001100110",
				"010001100110",
				"010001010101",
				"010001010101",
				"010001010101",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001010101",
				"011001100110",
				"011001110110",
				"011101110111",
				"100010001000",
				"100010011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101011001100",
				"101011001100",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101111101111",
				"101011101111",
				"101011101111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011001110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100011001101",
				"100011001101",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"100011001101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100011011101",
				"011111001100",
				"011110111100",
				"011110111100",
				"100011001101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011101",
				"011111001101",
				"100011001101",
				"100111011110",
				"100111001110",
				"100010111101",
				"011110111100",
				"011111001100",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111001101",
				"011110101011",
				"011010011010",
				"100010111011",
				"100111011101",
				"100011011101",
				"011011001100",
				"011111001100",
				"100110111101",
				"100010101100",
				"010101111001",
				"011110101011",
				"011111011101",
				"010111001100",
				"011111001100",
				"100011001101",
				"101011001101",
				"011110001010",
				"010001111000",
				"011010101011",
				"011111001101",
				"100011011101",
				"100111001101",
				"101010111100",
				"100110111011",
				"101010111100",
				"101111001110",
				"110011011111",
				"100110101101",
				"100010101101",
				"100110111110",
				"100010111110",
				"100010111101",
				"011110111100",
				"011010111011",
				"010111001100",
				"010111001100",
				"011011001101",
				"011111001101",
				"011111001101",
				"100010111110",
				"100011001110",
				"100011011110",
				"011110111100",
				"100010111011",
				"100110111011",
				"010101010101",
				"011001100110",
				"100010101010",
				"011110101010",
				"010110111011",
				"010111001100",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010101101",
				"011010111101",
				"010111001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011011001100",
				"010110111010",
				"011010111011",
				"011110111011",
				"011111001100",
				"011110111011",
				"011110111011",
				"011110111011",
				"100110111100",
				"100010101011",
				"011101111000",
				"100001111000",
				"011101111000",
				"011001100111",
				"100010011010",
				"100010101011",
				"011110111011",
				"011110111100",
				"011110111100",
				"011010101100",
				"010110101011",
				"010110111011",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110101011",
				"010110101010",
				"010010011010",
				"010010011010",
				"010110101010",
				"011010111011",
				"010110011001",
				"011110111011",
				"100011001011",
				"100010111011",
				"100011001100",
				"100011001100",
				"011010101010",
				"010001110111",
				"001101100111",
				"010001100111",
				"010101111000",
				"010110001001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101011",
				"011110101010",
				"011110011010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010101010",
				"011110111011",
				"010110011001",
				"010010001000",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001111000",
				"010110001000",
				"011010001001",
				"010101110111",
				"001101010101",
				"001001000101",
				"010001010110",
				"010001100111",
				"010001111000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110000111",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"010101111000",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010101111000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010101110110",
				"010101110111",
				"011001110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010101110110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001010101",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"001000110011",
				"010001000100",
				"010101010101",
				"011001100111",
				"011101110111",
				"100010001000",
				"100010001001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101110111100",
				"101011001100",
				"101011001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011111",
				"101011011111",
				"101111101111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011001110",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011101111",
				"101011011111",
				"101011101111",
				"101111011111",
				"101111101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"100011001101",
				"011110111101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011101",
				"100111011110",
				"100111011110",
				"100011011101",
				"100011001101",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011101",
				"100011001101",
				"011110111100",
				"011010101011",
				"011110111011",
				"100011001101",
				"100111011110",
				"101011011111",
				"100111011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011110",
				"100011001101",
				"011110111100",
				"011010111011",
				"011111001100",
				"100111011110",
				"100111011101",
				"100011001101",
				"100111001101",
				"100111011101",
				"100010111100",
				"100010111011",
				"100111001101",
				"100111011110",
				"100011011101",
				"011111001100",
				"100011001101",
				"100111001101",
				"100010101100",
				"011010011010",
				"100011001101",
				"011011001101",
				"010111001100",
				"011011001100",
				"100011001100",
				"101011001101",
				"011110011010",
				"001101100111",
				"011010011010",
				"100111011101",
				"101011011110",
				"100110111100",
				"100010101011",
				"100010111100",
				"101111101111",
				"101111011111",
				"101111011111",
				"100110111110",
				"100010101101",
				"011110101101",
				"100011001110",
				"100011001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011110111101",
				"011110111101",
				"100011001110",
				"011111001101",
				"011010111100",
				"011110111100",
				"101011001101",
				"101010111100",
				"011101100111",
				"011001100111",
				"100110101011",
				"011110111011",
				"011011001100",
				"011011001100",
				"010110111100",
				"010110111100",
				"011010111101",
				"011110111101",
				"010110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111101",
				"011110101100",
				"011010101100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"010110111011",
				"010110111011",
				"011010111011",
				"100010111100",
				"100010111100",
				"100010101011",
				"100110101011",
				"011101111000",
				"011101111000",
				"100010001001",
				"100110011011",
				"100010011010",
				"100110111100",
				"100011001101",
				"011110111011",
				"011010101100",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010011010",
				"010010011001",
				"010010011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011110011010",
				"100010101010",
				"010101111000",
				"010001100110",
				"010101110111",
				"010001110111",
				"001101100110",
				"001101010110",
				"010001110111",
				"011010001001",
				"011010011010",
				"011110011011",
				"011110101011",
				"011110101011",
				"011010101010",
				"011010101010",
				"010110011010",
				"011010101010",
				"010110001001",
				"010110011001",
				"011010011010",
				"011010101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"010110011001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110001001",
				"011010001001",
				"011010011001",
				"011010001000",
				"010101110111",
				"010101111000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"001110001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010101110111",
				"010001100110",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101100111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"001101010101",
				"010001100101",
				"010001100110",
				"010001100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001000110011",
				"010001000100",
				"010101010101",
				"011001100111",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101111011110",
				"101011011110",
				"101011011111",
				"101111101111",
				"101111101111",
				"101011011111",
				"101011011111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011001101",
				"100111001101",
				"101011001110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101011101110",
				"101011101110",
				"101011011110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011001110",
				"100111001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011110111101",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011101",
				"100111011101",
				"100111001101",
				"100111011101",
				"100011011101",
				"100011001101",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011101",
				"100111011101",
				"100111001101",
				"100111001101",
				"100111011110",
				"100111001101",
				"100111001101",
				"100011001101",
				"100010111100",
				"011110111011",
				"011110111100",
				"100011001101",
				"101011011110",
				"100111011110",
				"100111011110",
				"100011001101",
				"011110111100",
				"011111001101",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111001110",
				"100011001101",
				"011110111100",
				"100011001101",
				"100111011110",
				"100111011101",
				"100011001100",
				"100011001101",
				"100111011101",
				"100011001101",
				"100010111100",
				"100111001101",
				"100111011110",
				"100011011101",
				"100011011101",
				"100111011110",
				"101011001110",
				"100010101011",
				"011110101011",
				"100011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"100111011101",
				"100010101011",
				"010001100111",
				"011110011010",
				"101011001101",
				"100110111100",
				"011110011010",
				"100010101100",
				"100011001101",
				"100011001101",
				"100011001101",
				"101011101111",
				"101011011111",
				"011110101101",
				"011010101100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"100111011110",
				"101010111100",
				"011101111000",
				"010101000110",
				"100001111001",
				"100110101011",
				"011110111100",
				"011011001100",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"100010111101",
				"011110111101",
				"011010111100",
				"011010101011",
				"011110111100",
				"100011001100",
				"100011001100",
				"011111001100",
				"011111001100",
				"100011011101",
				"100011011101",
				"100011001101",
				"011110101011",
				"011010001001",
				"011110001010",
				"100010011011",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011110",
				"100110111100",
				"100111001101",
				"011110111100",
				"010110101011",
				"011010101011",
				"011010101100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010101011",
				"010110111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010001001",
				"011010001001",
				"011110011001",
				"011110001001",
				"010101100111",
				"001101000101",
				"001101000100",
				"010001100111",
				"011010001001",
				"011110011010",
				"011110011011",
				"011110011011",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010010011001",
				"010110011010",
				"011010101010",
				"010110011001",
				"011010101010",
				"011110101011",
				"011010101010",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"011010001001",
				"011110101010",
				"011010001000",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001111000",
				"010010001000",
				"010010011001",
				"010010001000",
				"001110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"001101100110",
				"001001010101",
				"001101010110",
				"010001110111",
				"010110001000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010001110111",
				"010001111000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110110",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101100110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"001000110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101111000",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111011110",
				"101111011110",
				"101011011110",
				"100111001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011001101",
				"100111011101",
				"100111011110",
				"100111011101",
				"100011001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"100011001101",
				"100111011110",
				"100111011101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100011001101",
				"100011001101",
				"100111001101",
				"100111011110",
				"101011101111",
				"100111011110",
				"100011001101",
				"011110111100",
				"011010101011",
				"011111001101",
				"100011011110",
				"100111101111",
				"100111011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"100011011101",
				"101011011110",
				"101011011110",
				"100011001100",
				"100011001100",
				"100111011110",
				"100011001101",
				"011110101011",
				"100111011101",
				"100111101110",
				"100011011101",
				"100111011110",
				"101011011110",
				"101111001110",
				"011110011010",
				"100010111100",
				"100011001101",
				"011111001101",
				"011011001100",
				"011111001101",
				"011111001100",
				"100011001100",
				"100010111011",
				"010001100111",
				"010101100111",
				"100010011010",
				"100010011011",
				"100010101011",
				"100010111101",
				"100011001101",
				"100011011110",
				"011111011101",
				"100011101110",
				"101011101111",
				"011110111100",
				"010010001010",
				"011110111100",
				"011111001101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"100011011101",
				"100011001101",
				"100010111100",
				"011110001001",
				"010101000110",
				"011101101000",
				"100110011011",
				"100110101100",
				"100010111101",
				"011110111101",
				"011010111101",
				"011111001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011110111100",
				"011010111100",
				"011110111100",
				"100010111100",
				"011010101011",
				"100010111011",
				"101011011101",
				"100110111100",
				"100010101011",
				"011110011010",
				"011010001010",
				"011010001010",
				"011010001010",
				"011110001010",
				"100010101100",
				"101011001101",
				"100110111101",
				"100010111100",
				"100010111100",
				"100011001100",
				"100011001101",
				"100111011101",
				"100011001101",
				"011110111100",
				"011010101100",
				"011010101100",
				"011010101011",
				"011010111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111100",
				"011010101011",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010011001",
				"011010011001",
				"011110011001",
				"011001110111",
				"001101000101",
				"010001010101",
				"011110001001",
				"100110011010",
				"100010011010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010011001",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010010011001",
				"010110101010",
				"010110011010",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011110101001",
				"011110011001",
				"010110001000",
				"010001100110",
				"001101010101",
				"010001010110",
				"010101110111",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"011010011001",
				"011010001000",
				"011010011000",
				"011110011001",
				"011010001000",
				"011010011000",
				"010110001000",
				"010110000111",
				"010001110111",
				"001101100110",
				"001001010101",
				"001101100110",
				"010001110111",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110110",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110110",
				"010001100110",
				"001101010101",
				"001101010101",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010010",
				"001000100011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"110011011111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100011011110",
				"100011001101",
				"100011001101",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"101011011110",
				"100111011110",
				"100011001101",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001101",
				"100011001101",
				"100011011101",
				"100111011110",
				"100111011101",
				"100111011110",
				"100111011110",
				"100111001101",
				"100011001101",
				"100011001100",
				"100011001101",
				"100111001101",
				"100111001101",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001101",
				"011110111100",
				"011010101011",
				"011110101100",
				"100011001110",
				"100111011110",
				"100111101110",
				"100111101110",
				"100011011110",
				"100011011110",
				"100011011101",
				"100111011110",
				"101011011110",
				"100111001101",
				"100010111100",
				"100011001101",
				"100111101110",
				"100111011101",
				"100011001100",
				"100111011110",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011001110",
				"100010011011",
				"011010001001",
				"100010111100",
				"100011001101",
				"011111001101",
				"011010111100",
				"011111001100",
				"011011001100",
				"011111001100",
				"100111011101",
				"011010001000",
				"010000110101",
				"011001010111",
				"100110011011",
				"100110111101",
				"100011001101",
				"100011001110",
				"011111011110",
				"011111101111",
				"011011011110",
				"100011101110",
				"100011011101",
				"010110011010",
				"010110011011",
				"011110111101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001100",
				"100011001101",
				"100111011101",
				"011110111011",
				"010101111000",
				"010001000110",
				"010101010111",
				"100110001010",
				"101010101101",
				"100110111101",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011010111100",
				"011111001100",
				"011110111100",
				"011010001001",
				"010101110111",
				"010101110111",
				"011001111000",
				"011001101000",
				"011110001010",
				"100010011011",
				"100010101100",
				"100010101101",
				"100110111101",
				"100010111101",
				"100010111101",
				"011110111100",
				"011111001100",
				"011111001100",
				"011010111011",
				"011010111011",
				"011110111100",
				"100010111101",
				"100011001101",
				"011110111100",
				"011010101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110011001",
				"011110011001",
				"011110001000",
				"010101100110",
				"100010001001",
				"100110011010",
				"100110101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010010101010",
				"010010101010",
				"010010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010110011010",
				"011010101010",
				"010110011010",
				"010010001001",
				"010110011001",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010101110111",
				"010001100110",
				"001101100101",
				"001101010101",
				"010001010101",
				"010101100110",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010110001000",
				"010110001000",
				"011010001000",
				"010101110111",
				"001101100110",
				"001001010101",
				"001001010101",
				"001001010101",
				"001101100110",
				"001101100110",
				"010001110111",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001100110",
				"010001110110",
				"010001110110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010001100111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011111",
				"101111011111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111001110",
				"100111011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100011001100",
				"011010111011",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100011001100",
				"100010111100",
				"100011001100",
				"100111001101",
				"100111001101",
				"100111001110",
				"100111001110",
				"101011011110",
				"100111001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111101111",
				"100011011101",
				"100011011110",
				"100011011110",
				"100111011110",
				"101011001101",
				"100010111100",
				"011110111100",
				"100011011101",
				"100111101110",
				"100011001101",
				"100010111100",
				"100111011110",
				"100111101111",
				"100111101111",
				"101011011110",
				"100110111100",
				"011010001001",
				"011010011010",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001100",
				"011111001011",
				"100111011101",
				"100110011010",
				"010101010110",
				"011101010111",
				"100110011011",
				"100010111100",
				"011111001101",
				"100011001111",
				"100011011111",
				"011111101111",
				"011011011101",
				"011011011101",
				"100011101110",
				"011110101100",
				"010001111001",
				"011010101100",
				"011110111110",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"100111011110",
				"100111011101",
				"101011001101",
				"100010101011",
				"010101111000",
				"010101111000",
				"011101111001",
				"011110001010",
				"100010011011",
				"011110011100",
				"011111001110",
				"011111001110",
				"011011001110",
				"011011001110",
				"011111001101",
				"011110111101",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011010111100",
				"011111001100",
				"100010111100",
				"011110101010",
				"010101100111",
				"010001000101",
				"011101101000",
				"100110001010",
				"101110101101",
				"101111001110",
				"100111001110",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011110111100",
				"100011001101",
				"011110111100",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110101011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010111011",
				"010110111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101001",
				"011110111010",
				"100110111011",
				"100010101010",
				"010001010110",
				"011110001001",
				"100010001010",
				"100010011010",
				"011010101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010101010",
				"010010011010",
				"010010011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011001",
				"010110011010",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011010011001",
				"011010011001",
				"011010001000",
				"011010001000",
				"011010011000",
				"011010011001",
				"011110011001",
				"011110011001",
				"011110001001",
				"011001110111",
				"010101100111",
				"010001100110",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"011010001000",
				"011010001000",
				"010101110111",
				"001101010101",
				"000100110100",
				"001101010101",
				"010001100110",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010110001000",
				"010001110111",
				"010001110111",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110000111",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001100110",
				"010001110110",
				"010101110111",
				"010101110111",
				"010001100111",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"001100110011",
				"010101010101",
				"010101010101",
				"011001100110",
				"011101110110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"101111011110",
				"101011001110",
				"101011001110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011001110",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011011111",
				"101011011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101111",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"101011011110",
				"101111011110",
				"100111011110",
				"011110111100",
				"011010111011",
				"011111001100",
				"100011011101",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100010111100",
				"011110111100",
				"011110111100",
				"100011001101",
				"100111011110",
				"101011011110",
				"101011011110",
				"100111001110",
				"100111001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"100011001101",
				"101011011111",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100011011110",
				"011111001101",
				"011111001101",
				"100011011110",
				"100111011110",
				"101011001101",
				"100010101100",
				"100010111100",
				"100111011110",
				"101011101111",
				"011110111100",
				"100010111100",
				"101011101111",
				"100111111111",
				"100011011110",
				"100111001110",
				"100110111101",
				"100010011011",
				"011110101011",
				"100011011101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100011011101",
				"011111001100",
				"100011011100",
				"100111011101",
				"100110101011",
				"011001010111",
				"011101101000",
				"100110011011",
				"011110111101",
				"100011011111",
				"100011001111",
				"100011011111",
				"011011001110",
				"011011011101",
				"011011011101",
				"011111011101",
				"100111011110",
				"010101111001",
				"011010001010",
				"100010111101",
				"011111001110",
				"011111011110",
				"100011011110",
				"100011001101",
				"100111011110",
				"100111001100",
				"011110011010",
				"100010101011",
				"100110111100",
				"101111001110",
				"100110111101",
				"011110001010",
				"011110011011",
				"011110111101",
				"011111001110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"010110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"011110001001",
				"010101010110",
				"100110001001",
				"110110111110",
				"101110101101",
				"100010101100",
				"011110101100",
				"011010111100",
				"010110111100",
				"010110111101",
				"011011001101",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010101100",
				"100010111101",
				"011110111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"010110101011",
				"010110101010",
				"011010101011",
				"011110111011",
				"100010111011",
				"100010101010",
				"011110011001",
				"010101100111",
				"010001010110",
				"011110001001",
				"100010011010",
				"011110011010",
				"011010101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110011001",
				"011010101010",
				"011110111011",
				"011110101011",
				"011010011010",
				"011010011010",
				"100010111011",
				"011110101011",
				"011110011010",
				"011010011001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010110001000",
				"011010001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"100010011010",
				"011110011001",
				"011110001001",
				"011010001000",
				"011010001000",
				"010110001000",
				"010010001000",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010110001000",
				"011010011000",
				"010110001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010101110111",
				"011010011001",
				"010110001000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010000111",
				"010010001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110110",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101100101",
				"011001100110",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011001101",
				"101011001101",
				"101111011101",
				"101111011110",
				"101111101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011111",
				"101011011111",
				"101011011111",
				"101111011110",
				"101011011110",
				"101011001110",
				"101011001101",
				"100111001101",
				"101011001110",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011101",
				"100011011110",
				"100111011110",
				"101111101111",
				"101111011110",
				"100111011110",
				"100010111100",
				"011111001100",
				"100011011101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100010111100",
				"011010101011",
				"011110111100",
				"100011001101",
				"100011011101",
				"100111011110",
				"101011011110",
				"101011011110",
				"100111001110",
				"100010111101",
				"011110111100",
				"011110111100",
				"100011001101",
				"100111011110",
				"101011011110",
				"100111001101",
				"101011011110",
				"101011011110",
				"100111011110",
				"011110111100",
				"011110111100",
				"011111001101",
				"100111011110",
				"101011101111",
				"101011001110",
				"100010111100",
				"100011001101",
				"100111011110",
				"100111011110",
				"011110111100",
				"100111001101",
				"101111101111",
				"100111101111",
				"011111001101",
				"100111001110",
				"101111011111",
				"100010111100",
				"011110111011",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111011110",
				"100011011101",
				"100011011101",
				"011111001100",
				"101011011101",
				"101010101011",
				"011001010110",
				"011001101000",
				"100110111101",
				"100011001110",
				"100011011111",
				"100011011111",
				"100011011111",
				"010111001101",
				"011011011110",
				"011011001101",
				"011111001101",
				"101011011110",
				"011110011011",
				"010101111001",
				"100010111100",
				"100111011110",
				"100111101111",
				"100111001110",
				"100010111100",
				"011110111100",
				"011110101011",
				"100010111100",
				"100111001101",
				"100111001101",
				"101011011110",
				"101111011111",
				"101111011111",
				"100111001110",
				"011010011011",
				"011010111101",
				"011111001110",
				"011111011111",
				"011011001110",
				"011011001101",
				"011111001101",
				"011011001101",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011011001101",
				"011111001101",
				"011110111100",
				"100110111100",
				"100110101011",
				"011001100111",
				"100010001001",
				"101010101100",
				"100010101100",
				"011010101100",
				"010110101100",
				"010110111101",
				"010111001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"011010101011",
				"011110101100",
				"100010111100",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010111100",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011110101011",
				"100010111100",
				"100010111100",
				"100010101011",
				"100010011010",
				"011101111000",
				"010001000101",
				"001100110100",
				"001101000101",
				"011110001001",
				"011110011010",
				"011110011010",
				"011110101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110011001",
				"011010011001",
				"011010011010",
				"011110101010",
				"011110101010",
				"011110011010",
				"011110011010",
				"010110001001",
				"010110001001",
				"010101111000",
				"010101111000",
				"010101111000",
				"010110001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011000",
				"010010001000",
				"001110001000",
				"001110001000",
				"001110001000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010011001",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010000111",
				"010110001000",
				"010110001000",
				"011110011001",
				"011110011001",
				"010110001000",
				"010110000111",
				"010101110111",
				"010110001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010001000",
				"010010000111",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"001101100110",
				"001101100110",
				"010001100110",
				"010001100110",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001100110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011001110111",
				"011110001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"101111001011",
				"101111001011",
				"101111001011",
				"101111001100",
				"101111001100",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101011001110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101011011111",
				"101111011111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011001110",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011011110",
				"100111001110",
				"100111011110",
				"101011011110",
				"101011101110",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011101110",
				"100111101110",
				"101111101111",
				"101111101111",
				"101011011110",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011101110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001101",
				"011110111100",
				"011010101011",
				"011110111100",
				"100111011110",
				"100011011110",
				"100111011110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100010111100",
				"011110111100",
				"100011001101",
				"100111101110",
				"100111011110",
				"101011011110",
				"101011001110",
				"101011011111",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111011110",
				"100111101111",
				"101011101111",
				"100111001110",
				"100111001101",
				"100011011110",
				"100011101110",
				"100111011110",
				"100011001101",
				"101011001110",
				"101011011111",
				"011111001101",
				"011011001100",
				"100111001101",
				"101111101111",
				"100010111011",
				"011110101011",
				"100011101110",
				"100011101111",
				"100111101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011101",
				"101011001100",
				"100110011010",
				"011001010111",
				"011001111001",
				"100111001101",
				"100011011111",
				"011111001110",
				"100011011111",
				"011010111101",
				"011011001110",
				"011011001101",
				"011011001101",
				"100011001101",
				"100110111101",
				"100110111101",
				"010101111000",
				"011010011010",
				"100010111100",
				"100111001101",
				"100010101100",
				"100010101011",
				"100010101100",
				"100010111100",
				"100010111101",
				"100111001110",
				"100011011101",
				"011111001101",
				"100011011110",
				"101011101111",
				"101111101111",
				"100111001110",
				"010110011011",
				"011010111101",
				"011111011110",
				"011111011111",
				"011011001110",
				"011011001101",
				"011011001101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011110111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011110111100",
				"101011001101",
				"101011001100",
				"100010001001",
				"011110001001",
				"011110001010",
				"100010111100",
				"100011001110",
				"011011001101",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111100",
				"011010101011",
				"011010101011",
				"011110101011",
				"011111001100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110011010",
				"011010001001",
				"011001111000",
				"010101100111",
				"010101010110",
				"010001010101",
				"010101010110",
				"010101010110",
				"100010101011",
				"011110011010",
				"011010011010",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010001001",
				"010110001000",
				"010110011001",
				"011010011001",
				"010110001000",
				"010001100111",
				"010001100111",
				"011010001000",
				"011110001001",
				"010101111000",
				"010101111001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010011000",
				"010010001000",
				"010010000111",
				"011010011000",
				"011110011001",
				"011110011001",
				"010101110111",
				"001101010101",
				"010001100110",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010010001000",
				"010010000111",
				"010010000111",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010101110111",
				"010001100110",
				"010001100110",
				"001101100110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101111000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010001110110",
				"010001100110",
				"010001100110",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100100010",
				"001000100010",
				"001101000100",
				"010001010101",
				"011001100110",
				"011001110111",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"101111011111",
				"101111011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101011001110",
				"101011001110",
				"101011001110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111101110",
				"101111101111",
				"101111011110",
				"101011011110",
				"100111011110",
				"100011011110",
				"100111101110",
				"100111101110",
				"100011011110",
				"100111011110",
				"100111011111",
				"100111011110",
				"100111001110",
				"100010111100",
				"011110111100",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"100010101100",
				"011110101100",
				"100010111101",
				"100111011110",
				"100111101110",
				"100111011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"100010111100",
				"100011001101",
				"100111101110",
				"101011011110",
				"101011011110",
				"100111101111",
				"100111011110",
				"100111001101",
				"100011001101",
				"100011101110",
				"100011101110",
				"101011101111",
				"100111001101",
				"101010111101",
				"100110111101",
				"011111001101",
				"011111011110",
				"100111011110",
				"101111101111",
				"100010111011",
				"011010101011",
				"100011101110",
				"100011111111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101110",
				"101011101110",
				"100110111011",
				"011001100111",
				"011001100111",
				"011110011010",
				"100011001101",
				"100011011111",
				"100011101111",
				"100011011110",
				"011011001101",
				"011011011110",
				"011011001110",
				"011110111101",
				"100010111110",
				"100010111101",
				"101011001110",
				"010110001001",
				"010001100111",
				"011110001001",
				"100010011010",
				"100010001010",
				"100110101100",
				"100110111101",
				"100111001110",
				"011110111101",
				"011111001110",
				"011011011101",
				"011011101110",
				"011111011101",
				"011111001101",
				"101011011110",
				"101111011111",
				"011110101100",
				"010110101011",
				"011010111100",
				"011111011110",
				"011111011110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011110111100",
				"100110111100",
				"100110101011",
				"100010001001",
				"011110001001",
				"011110011011",
				"011110111100",
				"011111001101",
				"011010111101",
				"010111001101",
				"011011001110",
				"011011001101",
				"011010101100",
				"011010101100",
				"011010101011",
				"010110101010",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"011110111011",
				"011010101011",
				"011010101011",
				"011110111100",
				"100011001101",
				"011111001101",
				"011110111100",
				"011010101011",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100011001100",
				"100011001100",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010101011",
				"011110011011",
				"010110001001",
				"010001111000",
				"001101100111",
				"010001111000",
				"010110001001",
				"100010101011",
				"100110111100",
				"100110111100",
				"011110011001",
				"011110101010",
				"011010011010",
				"011010011010",
				"011010011011",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"010101110111",
				"010001010110",
				"010101110111",
				"011110001001",
				"011010001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"001110001000",
				"010010011001",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011110101010",
				"011010001000",
				"011001110111",
				"010001010110",
				"010001010101",
				"010001010110",
				"010101100110",
				"010101110111",
				"010101110111",
				"010110001000",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110000111",
				"010110001000",
				"010110000111",
				"010110000111",
				"010110000111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110110",
				"010101110111",
				"010101110111",
				"010101111000",
				"010101110111",
				"010101110111",
				"010101100111",
				"010101110111",
				"010101111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101111000",
				"010101111000",
				"010101110111",
				"010101111000",
				"010101111000",
				"010001110111",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110000111",
				"010110001000",
				"010110000111",
				"010001110111",
				"010001100110",
				"001101100110",
				"001101010101",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001101000100",
				"010001010101",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"101111001100",
				"101111001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"101111011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011011111",
				"110011011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111001110",
				"101011001110",
				"101011001110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101111011110",
				"101111101111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111101111",
				"101111011111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011011110",
				"100111011110",
				"100111101110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111101111",
				"100111101111",
				"100111011110",
				"100111011110",
				"101011011111",
				"100111011110",
				"100111011110",
				"100111001101",
				"100011001101",
				"100011011110",
				"100111101110",
				"100111101110",
				"100111001101",
				"100010101100",
				"011010011011",
				"011110101100",
				"100011001101",
				"100111101111",
				"100111101111",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111001101",
				"100010111100",
				"100111011101",
				"100111011110",
				"101011011111",
				"101011011111",
				"101011101111",
				"100111011110",
				"100010111100",
				"100011001101",
				"100011101110",
				"100011101110",
				"101011101110",
				"011110101011",
				"011110001010",
				"011110001010",
				"011111001101",
				"100111101111",
				"100111011110",
				"101011101111",
				"011110111100",
				"011010111011",
				"100011101110",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011111111",
				"100111011110",
				"100010111011",
				"011110001001",
				"010101010110",
				"011101111001",
				"100110111101",
				"100011011110",
				"100011101111",
				"011111011111",
				"011111011110",
				"100011101110",
				"011111011110",
				"011111011110",
				"100011001110",
				"100010111110",
				"100010111101",
				"100111001101",
				"100010101011",
				"010001100110",
				"011101111000",
				"100110001001",
				"100110011011",
				"101110111110",
				"100110111110",
				"100011001110",
				"100011011111",
				"011111011110",
				"010111011110",
				"011011101110",
				"011011101110",
				"011011001101",
				"100011001101",
				"100111001101",
				"100111011110",
				"011010101011",
				"010010101011",
				"011011001101",
				"011111011110",
				"011011001110",
				"011011001110",
				"011111001110",
				"011011001101",
				"011011001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100111001110",
				"101011001110",
				"100010101011",
				"011001111000",
				"011110001001",
				"100110101011",
				"100010101100",
				"011110111100",
				"011110111101",
				"011011001101",
				"010110111100",
				"010110111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101010",
				"010010101010",
				"010010101010",
				"010110111011",
				"011010111100",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011110111100",
				"100011001101",
				"011110111100",
				"011110101100",
				"100010111100",
				"100110111101",
				"100110111100",
				"100010111100",
				"011110101011",
				"011010101010",
				"010110011001",
				"011010001001",
				"011001111001",
				"010101111001",
				"011010011010",
				"011010011010",
				"010110101010",
				"011010101011",
				"011111001100",
				"011110111100",
				"011110111011",
				"100011001100",
				"100011001100",
				"100010111100",
				"100010111100",
				"011110011011",
				"010110001010",
				"011010011010",
				"011010101011",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110011001",
				"011010001000",
				"011010001000",
				"011110011001",
				"011110011010",
				"011110101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110001000",
				"010001100110",
				"001101010101",
				"001000110100",
				"001101000101",
				"010101100110",
				"010001010110",
				"010001100110",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010110001000",
				"010010001000",
				"010010000111",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010110000111",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110000111",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"010101110111",
				"010101110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010101111000",
				"010101111000",
				"010101111000",
				"010001110111",
				"010010000111",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001100111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011001100",
				"110111001100",
				"110111001101",
				"110111011101",
				"110011011100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011011111",
				"101111011110",
				"101111001110",
				"101111001101",
				"101011001101",
				"101111011110",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101011001101",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101110",
				"101111101110",
				"101111101110",
				"110011101111",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111011110",
				"101011001110",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011101110",
				"101111101110",
				"101111101110",
				"101111101110",
				"101011011110",
				"100111011110",
				"101011101110",
				"100111101110",
				"100111101110",
				"100111101110",
				"100111011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111011110",
				"100111001101",
				"011110011010",
				"011010011010",
				"100010111101",
				"100111101111",
				"100011011110",
				"101011101111",
				"101011011111",
				"100111001101",
				"100010111100",
				"100010111100",
				"100011001101",
				"101011011110",
				"100111011101",
				"100111011110",
				"101111111111",
				"101111011110",
				"100010101011",
				"100010111100",
				"100111011101",
				"100011101110",
				"100011101110",
				"100111011110",
				"011110101011",
				"001101010111",
				"011110011011",
				"100111001110",
				"100111101111",
				"100011011110",
				"100111101111",
				"011111001101",
				"011011001100",
				"100011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"100011001101",
				"100010001010",
				"011101101000",
				"011101111001",
				"100110101100",
				"100110111101",
				"100011011110",
				"011111011111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100011101111",
				"011111011110",
				"011011011110",
				"011011011110",
				"011111011101",
				"011111001100",
				"100111001100",
				"011010001000",
				"011001100111",
				"100010001001",
				"101110111100",
				"101010111110",
				"011110111101",
				"011111011111",
				"011111001110",
				"011111001110",
				"011011011110",
				"011011011110",
				"011011011101",
				"011011001101",
				"011111001101",
				"100011001101",
				"100011011110",
				"100111011110",
				"010110101011",
				"010110101011",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001111",
				"011111011111",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111001101",
				"011110111100",
				"100111001100",
				"101111001101",
				"101010101011",
				"100001111000",
				"011001100111",
				"100010001010",
				"101010111100",
				"101011001101",
				"011110101100",
				"100011001110",
				"011110111101",
				"010110111100",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111100",
				"100010111100",
				"011010001001",
				"011110001010",
				"100001111001",
				"011001010111",
				"011001101000",
				"011110001001",
				"010110001000",
				"011010011001",
				"100010101011",
				"100010101100",
				"011110101100",
				"011110101011",
				"011010111100",
				"011011001100",
				"010111001100",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"100010111100",
				"100010101100",
				"011110101011",
				"011010011010",
				"010110011001",
				"010110011010",
				"011010011011",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010111011",
				"010010011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010011001",
				"011110011001",
				"011110011001",
				"011010001000",
				"100010101010",
				"010110001000",
				"011010001000",
				"011010011001",
				"011010011010",
				"011010101011",
				"011010101011",
				"010110011010",
				"010010011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011001",
				"010110001001",
				"010010001000",
				"010110011001",
				"010010001000",
				"010110011001",
				"010110011010",
				"011010101010",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010110001001",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010011001",
				"010001111000",
				"001101100110",
				"001101100110",
				"010001100111",
				"010101111000",
				"010110001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010001110111",
				"001101110111",
				"010010001000",
				"010110011000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011000",
				"010110001000",
				"010010000111",
				"010010000111",
				"010110001000",
				"010110001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"011010001000",
				"011010001000",
				"011010001001",
				"011010001001",
				"010101110111",
				"001101100110",
				"010001110111",
				"010010001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001110111",
				"010110001000",
				"011010011001",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101111000",
				"010101111000",
				"010101110111",
				"010001100110",
				"001101100110",
				"001101010101",
				"001101010101",
				"001101100110",
				"010001100110",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100110",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101011",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110111001100",
				"110111001100",
				"110111011100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001011",
				"110011001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011011110",
				"110011011110",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011110",
				"101111101110",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011011101",
				"101011011110",
				"101011101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011111",
				"101111101111",
				"101011101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101110",
				"101111101110",
				"101111101110",
				"101111101110",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111011110",
				"101011001110",
				"101011001110",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011101110",
				"101011101110",
				"101011101110",
				"101011101111",
				"101011101110",
				"101011101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111011110",
				"100110111101",
				"011110011011",
				"011110101011",
				"100011001101",
				"100111101110",
				"100111011110",
				"101011011111",
				"100111001101",
				"011110101100",
				"100010111100",
				"100011001101",
				"100111011101",
				"101011011110",
				"100111001101",
				"100111011110",
				"101011011110",
				"101011001101",
				"101010111101",
				"101011011101",
				"101011011110",
				"100011101110",
				"100011101110",
				"100111101110",
				"011110111100",
				"010001111000",
				"100010111100",
				"101011011111",
				"101011101111",
				"100011101111",
				"100111111111",
				"011111001101",
				"011110111100",
				"101011101111",
				"100111011110",
				"101111101111",
				"101011101111",
				"011111001100",
				"100111001101",
				"101110111101",
				"101110101100",
				"100010001010",
				"100110101100",
				"100111001101",
				"100111011111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011011011110",
				"011011011101",
				"011011011101",
				"100011011101",
				"101111011101",
				"100010011001",
				"011001100111",
				"100110011001",
				"101010111101",
				"100110111101",
				"011111001110",
				"011011011111",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011011001101",
				"011111001101",
				"011111011110",
				"100011011110",
				"011110111100",
				"010110011011",
				"011010111100",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"100011011110",
				"100011011101",
				"100111001101",
				"101011001101",
				"100110101010",
				"100010001001",
				"100010001001",
				"100110001010",
				"100110011010",
				"100110101100",
				"100111001101",
				"100011001110",
				"011010111101",
				"011010111101",
				"011111001110",
				"011010111101",
				"011010111101",
				"011111001101",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110101011",
				"100010101011",
				"011001111000",
				"011001010110",
				"011101100111",
				"100110001001",
				"100110101011",
				"100110111011",
				"011110101010",
				"011110101011",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010010111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011110111100",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010011010",
				"011010011010",
				"011010101011",
				"011110101100",
				"011010101011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010101010",
				"010110101010",
				"010110101001",
				"011010101010",
				"011010011001",
				"011010001001",
				"011110011001",
				"011110011001",
				"011110011001",
				"001101010110",
				"010001100110",
				"011010011010",
				"010110011010",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010001001",
				"011010011010",
				"100010111011",
				"011010011010",
				"011010011010",
				"010110001001",
				"001101100111",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110011000",
				"010110011000",
				"010110001000",
				"010110011000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110011000",
				"010110011000",
				"010110011000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011110011001",
				"011001111000",
				"011010001000",
				"011110001001",
				"010101100111",
				"010001100110",
				"010101110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010010001000",
				"010110001000",
				"010110001000",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001100111",
				"001101010101",
				"001101010101",
				"001101010101",
				"001101010110",
				"001101100110",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001110111",
				"001101110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011110000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110111001100",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001011",
				"101111001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"101111001110",
				"101111001101",
				"101111001101",
				"101111011110",
				"101111101110",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011001101",
				"101011011110",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111101110",
				"101111101110",
				"101111101110",
				"101111101110",
				"101111011110",
				"101111011110",
				"101111011111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101011011101",
				"100111011101",
				"101011011110",
				"101011101110",
				"101011101110",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"100111101110",
				"100111101110",
				"101011011110",
				"100111001101",
				"100010101100",
				"100010111101",
				"100111011110",
				"100111011110",
				"100111101111",
				"101011011110",
				"100010111100",
				"011010011010",
				"011110101100",
				"100111001101",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111011110",
				"100111001101",
				"100111001101",
				"101111011110",
				"101111101111",
				"101011101110",
				"100111011110",
				"100111101110",
				"101011101110",
				"100010111100",
				"010110001001",
				"100111001101",
				"101011101111",
				"100111101111",
				"100011011111",
				"101011111111",
				"011110111100",
				"100010111100",
				"101011011110",
				"101111101111",
				"101111101111",
				"011111001100",
				"011011001100",
				"100111101110",
				"110011101111",
				"110011001110",
				"100010011010",
				"100010011011",
				"100111001101",
				"100111011111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111011110",
				"011111001101",
				"100111001101",
				"110011101110",
				"100110011001",
				"011001100110",
				"100110011010",
				"100110111101",
				"011110111101",
				"011111011111",
				"011011011111",
				"011011011111",
				"011111011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111001110",
				"011011011101",
				"011011011101",
				"011011011101",
				"011111001101",
				"100011001110",
				"011010011011",
				"011010011011",
				"100010111101",
				"100011011110",
				"100011011110",
				"011111001101",
				"100011001110",
				"100011001110",
				"100111011111",
				"101011011111",
				"100111001110",
				"100010111100",
				"011110101011",
				"100010101011",
				"101011001100",
				"110011101110",
				"110011101111",
				"101111001110",
				"101010111101",
				"101010111101",
				"101011001110",
				"011110101100",
				"011111001101",
				"011111001110",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"011010101010",
				"100010111100",
				"100010101011",
				"011001111000",
				"011101111001",
				"100110101011",
				"100010011010",
				"011110101010",
				"011110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011110111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101011",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110111010",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010111011",
				"010110101010",
				"010010101001",
				"010010101010",
				"010110111010",
				"011010111011",
				"011010101010",
				"011010011010",
				"100010101011",
				"100010101011",
				"011110001001",
				"010001010110",
				"010101010110",
				"011001111000",
				"011001111000",
				"011110001001",
				"011010011011",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011110011010",
				"011110011010",
				"011110011010",
				"010001111000",
				"001101100110",
				"001101100110",
				"001101100110",
				"001101100110",
				"010001110111",
				"010001111000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010001111000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011000",
				"010010001000",
				"010110001000",
				"010110011000",
				"011010011001",
				"011110001001",
				"011110001000",
				"011001111000",
				"011001110111",
				"010101100111",
				"010001010110",
				"010001010110",
				"010001100111",
				"010001110111",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110000111",
				"010110000111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010101110111",
				"010001100111",
				"010001100110",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100111",
				"010001100111",
				"010001100111",
				"010001100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"110010111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"101111001011",
				"101111001011",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011111",
				"110011011110",
				"110011011110",
				"101111001101",
				"101111001101",
				"101111011110",
				"110011101110",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011011111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101011001101",
				"101011011101",
				"101011011110",
				"101111101111",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101011101110",
				"101011101110",
				"100111011110",
				"101011101110",
				"101011101110",
				"100111001101",
				"100110111100",
				"101011011110",
				"101011011110",
				"100111011110",
				"101011101111",
				"101011011110",
				"011110101011",
				"011010011010",
				"100010111100",
				"100111011110",
				"101011101110",
				"101011011110",
				"100111001101",
				"100111001101",
				"100010111100",
				"100111001101",
				"101111101110",
				"101011101110",
				"100111011110",
				"101011101110",
				"101111101111",
				"101011011110",
				"100010101011",
				"011010011010",
				"100111011110",
				"100111101111",
				"100011101111",
				"100011011111",
				"101011101111",
				"100010111100",
				"100010111100",
				"101111011110",
				"110011101111",
				"100111001101",
				"011010111100",
				"100011101110",
				"100011101110",
				"101011101111",
				"101111011110",
				"011110011010",
				"011010001010",
				"100011001101",
				"100111011111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111011111",
				"100111011110",
				"101011011110",
				"110011011101",
				"100010001001",
				"011101100111",
				"100110101010",
				"100011001101",
				"011111001101",
				"011111011111",
				"011111011111",
				"011011011111",
				"011011011110",
				"011111001110",
				"100010111110",
				"100010111110",
				"011111001110",
				"011011011110",
				"011011011110",
				"010111011101",
				"011011001101",
				"100111001110",
				"100010111100",
				"011110011010",
				"100010101100",
				"100011001101",
				"100111011110",
				"100111011110",
				"101011011111",
				"101011011111",
				"101011001110",
				"100110111101",
				"011110101011",
				"011110101011",
				"011110101100",
				"100011001101",
				"100111011101",
				"100111011101",
				"100111001101",
				"101011011110",
				"101111101111",
				"101011011111",
				"100010101100",
				"011010011011",
				"011110111101",
				"011111001110",
				"011110111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011110111011",
				"100010111100",
				"011110001001",
				"011001111001",
				"100110101011",
				"100010101011",
				"011010101010",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101010",
				"011110111011",
				"011110111100",
				"010110101011",
				"010010101010",
				"010110111011",
				"011010111100",
				"011010101011",
				"011110111100",
				"011010111011",
				"011010111011",
				"010110111010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110101010",
				"011010101010",
				"011110111011",
				"011010001001",
				"010001100111",
				"001101000101",
				"001000110100",
				"010001000101",
				"011101111001",
				"011001111000",
				"011110011010",
				"011110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"001101010110",
				"001001000101",
				"001101010110",
				"010001100111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001111000",
				"010110001000",
				"011010011010",
				"011010011001",
				"010110001000",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010001110111",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011000",
				"010110011001",
				"011010011001",
				"010110001000",
				"010001111000",
				"010001111000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011001111000",
				"011001111000",
				"011110001001",
				"010101110111",
				"010001010110",
				"010001100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010001110111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010101110111",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010101010100",
				"010101010101",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110111001100",
				"110111001100",
				"110011001100",
				"110011001011",
				"101110111011",
				"101110111011",
				"101111001011",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011101110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"101111001101",
				"101111011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101011001110",
				"100111001110",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111011111",
				"110011101111",
				"110011101111",
				"110011011111",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011001101",
				"101011011101",
				"101111101110",
				"101111101111",
				"101111101110",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111001110",
				"101011001101",
				"101111011110",
				"101111011111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101111101111",
				"101011011110",
				"100111001101",
				"100111001101",
				"101011011111",
				"101011101111",
				"100111011110",
				"101111101111",
				"101011011110",
				"011110101011",
				"011110101011",
				"100011001101",
				"101011101110",
				"101011101110",
				"100111001101",
				"100110111100",
				"100010101011",
				"100111001101",
				"101011011110",
				"101011011110",
				"100111011110",
				"101011101110",
				"101111101111",
				"101111101111",
				"101010111101",
				"011110011010",
				"011010101011",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101111101111",
				"100110111100",
				"100010011011",
				"101111001110",
				"100110111100",
				"011010101011",
				"100011011110",
				"100011101111",
				"100011011110",
				"101011101111",
				"101111101111",
				"011110101011",
				"010110001001",
				"011110111100",
				"100011011110",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101010101011",
				"011101111000",
				"100010001000",
				"100010101011",
				"011111001101",
				"011111011110",
				"011111011111",
				"011111101111",
				"011111011111",
				"011111011110",
				"011111001110",
				"100011001110",
				"100010111110",
				"011111001110",
				"011011001110",
				"011011011110",
				"011011011101",
				"011011001101",
				"100011001101",
				"100111001110",
				"100010101011",
				"011010001001",
				"100010101011",
				"100010111100",
				"100110111100",
				"100010111100",
				"100010101011",
				"100010101011",
				"100010101100",
				"100110101100",
				"100110111101",
				"100111001110",
				"100111011110",
				"100011011110",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011001110",
				"101011011111",
				"101011101111",
				"100011001110",
				"011010101011",
				"011110111100",
				"100011001110",
				"011110111100",
				"011010101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"011011001100",
				"011011001100",
				"011011001011",
				"011011001011",
				"011010101010",
				"011110101011",
				"100010101011",
				"011010001001",
				"011010001001",
				"100010101011",
				"011110111100",
				"010110101011",
				"010110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010011010",
				"011110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010101011",
				"011010101010",
				"011010111011",
				"011010111100",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101010",
				"010110101010",
				"011010111010",
				"100010111100",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"011010111011",
				"011010111011",
				"011010101010",
				"010110011001",
				"010001111000",
				"010001100111",
				"010101110111",
				"010101111000",
				"010101100111",
				"010101111000",
				"100010101011",
				"011010001000",
				"010101111000",
				"011010101010",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"011010101001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010101110111",
				"001001000101",
				"010001010110",
				"011001111000",
				"011010001001",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001000",
				"010110001000",
				"011010001000",
				"010101110111",
				"011010001000",
				"011110011001",
				"011010011001",
				"011010011001",
				"011010011001",
				"010101111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010001110111",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001100111",
				"011010001000",
				"010101110111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"110011001011",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011110",
				"110011011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011101111",
				"101111101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011111",
				"101111011111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011011101",
				"101011011110",
				"101111101110",
				"101111101111",
				"101111101110",
				"101111101110",
				"110011101111",
				"110011011110",
				"101111001101",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"100111001101",
				"101011001101",
				"101111101111",
				"101011101111",
				"101011011110",
				"101111101111",
				"101011011110",
				"100010111100",
				"100010111100",
				"100111011101",
				"101011101110",
				"100111011110",
				"100010111100",
				"100010101011",
				"100010101011",
				"101011001101",
				"101011101110",
				"100111011110",
				"100111101110",
				"101111111111",
				"101111101111",
				"101111001110",
				"100110101011",
				"011010001001",
				"011110111100",
				"100111101111",
				"100011111111",
				"100011101111",
				"100111101111",
				"101011101111",
				"100110111100",
				"011001111001",
				"011001111001",
				"011010001010",
				"100010111101",
				"100011011110",
				"100011101110",
				"100011101110",
				"100111101111",
				"101111111111",
				"100010111100",
				"010001111001",
				"011010101011",
				"100011011110",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101011001110",
				"100110101100",
				"100001111001",
				"011101101000",
				"100110011010",
				"100010111100",
				"011111011101",
				"011111101111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"011111001110",
				"011011001110",
				"011011001101",
				"011011011110",
				"011011001101",
				"011010111100",
				"100111011110",
				"100010111100",
				"010101111000",
				"011001111000",
				"011110001001",
				"011010001001",
				"011110001001",
				"011110011010",
				"100110101100",
				"101010111101",
				"101011001110",
				"100111001110",
				"100011001101",
				"100011001110",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"100011001110",
				"100111011111",
				"011110111100",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011010111100",
				"011111001101",
				"011011001101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001011",
				"011111001011",
				"011110111011",
				"100010111100",
				"100110111100",
				"011001111001",
				"010101111000",
				"011110101011",
				"011010101011",
				"010110101011",
				"010110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101010",
				"011110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010101010",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010011010",
				"011110101010",
				"011110101011",
				"100011001100",
				"100011001100",
				"011110111011",
				"100010111011",
				"100010111100",
				"100010111011",
				"100010111011",
				"011110101011",
				"011110101011",
				"010110001001",
				"001101110111",
				"001001010110",
				"001001100110",
				"001101100111",
				"011110101011",
				"011110101011",
				"100010111011",
				"100111001100",
				"100010111100",
				"100010111100",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"011001111000",
				"011001111000",
				"011001111000",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"011010001001",
				"011010001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"011010001000",
				"010110001000",
				"010110011000",
				"011010011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010010001000",
				"010010001000",
				"010010000111",
				"010001110111",
				"010010000111",
				"010010001000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010001000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010110001000",
				"010001110111",
				"010001100111",
				"010001100111",
				"010001110111",
				"010001111000",
				"010001110111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100011",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101111000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"110010111011",
				"110010111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"101011001101",
				"101011001110",
				"101011011110",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"101011001101",
				"101011011101",
				"101011011110",
				"101111101110",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101011011110",
				"101111011110",
				"101111101110",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111101110",
				"101111101110",
				"101111011110",
				"101111101110",
				"110011101111",
				"110011011110",
				"101111001101",
				"101010111101",
				"101011001101",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011001101",
				"100111001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101011011110",
				"100110111100",
				"100111001101",
				"100111011110",
				"101011101110",
				"101011011110",
				"100010101011",
				"011010001001",
				"100010101011",
				"101011011110",
				"101111101111",
				"100111011110",
				"101011101110",
				"101111101111",
				"101111011110",
				"101011001101",
				"100110101100",
				"011010001001",
				"100011001101",
				"101011111111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011011111",
				"101011001101",
				"010101101000",
				"001101000110",
				"011110011011",
				"101011101111",
				"100011011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"100111001101",
				"010001111000",
				"011010101011",
				"100011101110",
				"100011101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011011111",
				"101111101111",
				"101011101111",
				"100111011110",
				"011110101011",
				"011101111001",
				"100001111001",
				"101010011010",
				"101010111100",
				"100011001100",
				"011111011110",
				"011111101111",
				"011111101111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011111",
				"011111011110",
				"011111001110",
				"011011001110",
				"011011001110",
				"011011001101",
				"011011001100",
				"100011011101",
				"100111001101",
				"011110001001",
				"011001100111",
				"011101111000",
				"100110011010",
				"101010111100",
				"101111001101",
				"100111001101",
				"100010111100",
				"011110111100",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"100111011110",
				"011110111100",
				"010110011010",
				"011110111100",
				"100011001110",
				"011110111101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011111001100",
				"011110111100",
				"100010111011",
				"100010111011",
				"100010111011",
				"100010011010",
				"011001111001",
				"011001111001",
				"011110011011",
				"100010111100",
				"011010101100",
				"010110101100",
				"010110101100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101010",
				"011010101011",
				"011010101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110101011",
				"011010011010",
				"011110101010",
				"011110011010",
				"100110111011",
				"100110111011",
				"100010101010",
				"011110011001",
				"011110011001",
				"011010001001",
				"011001111001",
				"010101111000",
				"010001100111",
				"010001101000",
				"010101111000",
				"011010011010",
				"011110101011",
				"100010111100",
				"011010101010",
				"011110111011",
				"011110111011",
				"011010101010",
				"010110101010",
				"011111001100",
				"011111001100",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"010101111000",
				"011110001001",
				"011110011001",
				"011101111001",
				"010001010110",
				"011010001001",
				"011010011010",
				"010110001000",
				"010110011001",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011000",
				"010010011000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"011010011001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"011110011010",
				"011010001001",
				"010110001001",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"011010011001",
				"010110001000",
				"010001110111",
				"010010001000",
				"010010000111",
				"001101110111",
				"010110011000",
				"010110011001",
				"010110001001",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"001101010110",
				"001101010110",
				"001101010110",
				"001101100110",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101100111",
				"001101110111",
				"001101100111",
				"001101100111",
				"001101110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110111011101",
				"110011011101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"101011001110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101011101111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011001110",
				"100111001101",
				"101011001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111101110",
				"101111101110",
				"101111011110",
				"101111101110",
				"110011101111",
				"110011011110",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011110",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111001110",
				"101010111101",
				"100111001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"100111001101",
				"100111011110",
				"101011011110",
				"101011101111",
				"101011011110",
				"011110101011",
				"010101111000",
				"100010111100",
				"101011011110",
				"101111101111",
				"101011011110",
				"101011101110",
				"101011011110",
				"101011011110",
				"101111001110",
				"101010111101",
				"011110011011",
				"100111011110",
				"101011111111",
				"100011101110",
				"100011101111",
				"101011101111",
				"101011011111",
				"101111101111",
				"010001100111",
				"010101111001",
				"100010111100",
				"100111011110",
				"100111101111",
				"100111101111",
				"100011011110",
				"100111101111",
				"101011101111",
				"101011011110",
				"010101111000",
				"011010011010",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111101111",
				"110011101111",
				"101111101111",
				"100011011110",
				"011010111100",
				"011110101011",
				"100110101100",
				"100110001010",
				"110010111101",
				"101011001101",
				"100011001101",
				"011011011101",
				"011111101111",
				"100011111111",
				"011111011111",
				"011111101111",
				"011111101110",
				"011111011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"011011001110",
				"011011001101",
				"011011001101",
				"011111001101",
				"101011011110",
				"100110111100",
				"011101101000",
				"100001111000",
				"101010101011",
				"101010111100",
				"100110111100",
				"011110111100",
				"011110111101",
				"011111001110",
				"100011011110",
				"011111001110",
				"011111001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"011011001101",
				"011011001101",
				"011011001110",
				"011111011110",
				"011111011101",
				"100011011101",
				"011111001101",
				"011110111100",
				"011010111100",
				"011110111100",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011110111101",
				"011110111100",
				"100010111100",
				"100010111100",
				"100110111100",
				"100110111100",
				"100010011010",
				"011001101000",
				"011001101000",
				"100110101100",
				"100010101100",
				"011010011011",
				"011110111101",
				"011010101100",
				"010110101100",
				"011010111100",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111010",
				"011010111010",
				"011010111010",
				"011010111010",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"100010111100",
				"010110001000",
				"010001100110",
				"010101100110",
				"011001100111",
				"010101010110",
				"010001010110",
				"010101111000",
				"011010001000",
				"010101111000",
				"011001111001",
				"011010001010",
				"011110011011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010111011",
				"010110101011",
				"010010101010",
				"010110111011",
				"011011001100",
				"011111001100",
				"011010101010",
				"010010011001",
				"010110011001",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110101001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010101111000",
				"011010001001",
				"011110001001",
				"011110001001",
				"010101100111",
				"010001100111",
				"011010011010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001001",
				"011110001001",
				"010101111000",
				"010101111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010010000111",
				"010010001000",
				"001101110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"010001100111",
				"010101110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101110",
				"101111101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101111101110",
				"101011011110",
				"101011011101",
				"101111011110",
				"110011101110",
				"110011011110",
				"101111001110",
				"101011001101",
				"101111001101",
				"110011101110",
				"101111101111",
				"101111101110",
				"101011101110",
				"101111101110",
				"101111001101",
				"101011001101",
				"100111001101",
				"101011011110",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111011110",
				"101010111100",
				"100111001101",
				"101011011110",
				"101011101110",
				"101011101110",
				"101011011110",
				"011110011010",
				"011110011010",
				"100111001101",
				"101011011110",
				"101111101111",
				"101011011110",
				"101011011110",
				"100111001101",
				"101011001101",
				"110011101111",
				"101010111101",
				"100010101011",
				"101011011111",
				"100111101110",
				"100111101111",
				"100111111111",
				"100111101110",
				"101011101111",
				"101111101111",
				"011010001001",
				"010001101000",
				"100111001101",
				"100111011110",
				"100111101111",
				"100111101111",
				"100011101110",
				"100011101111",
				"101011111111",
				"101111101111",
				"011010001001",
				"010110001001",
				"101011011110",
				"100111011110",
				"101111111111",
				"101111101111",
				"110011111111",
				"110011011111",
				"100010101100",
				"010110101011",
				"011111011101",
				"101011101111",
				"101111011111",
				"101110111101",
				"101010101100",
				"101011001101",
				"011110111100",
				"011111011110",
				"011111101111",
				"011111101111",
				"100011101111",
				"011111101111",
				"011111101110",
				"011111011110",
				"100011011110",
				"100011011111",
				"100011011111",
				"011111011110",
				"011011001110",
				"011011011110",
				"011011001101",
				"011111001101",
				"100010111100",
				"101011011110",
				"101010111100",
				"011101100111",
				"100001111000",
				"101010101011",
				"100110111100",
				"100011001101",
				"011111001101",
				"011011011110",
				"011011011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"100011101110",
				"010110111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011011001101",
				"011111011101",
				"011111001101",
				"011110111100",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100110111100",
				"100010011011",
				"100010001010",
				"100001111001",
				"100001111001",
				"100110001011",
				"100110101100",
				"100010101100",
				"011110101100",
				"011111001110",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011110101010",
				"011010001000",
				"001100110100",
				"010001000101",
				"011001100111",
				"011001111000",
				"100010101011",
				"011110101011",
				"011010011010",
				"011110101011",
				"011010101011",
				"011010011010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"011010111011",
				"011110101011",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110101001",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011110011010",
				"011110011001",
				"010101110111",
				"010101010110",
				"010001010110",
				"010101111000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001100110",
				"001101010110",
				"010101100111",
				"011010001001",
				"010110001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010001110111",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010001110111",
				"001101100110",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100011",
				"010001000100",
				"010101010101",
				"011001010101",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001011",
				"110011001011",
				"110011001011",
				"101111001011",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011101110",
				"110011101110",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"110011011110",
				"110011101111",
				"110011011111",
				"110011101111",
				"101111101111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011101",
				"101111011110",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011011110",
				"101011011110",
				"101111101110",
				"101111001101",
				"101111001101",
				"101011001101",
				"101111101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111001101",
				"100110111100",
				"100111001101",
				"101011011110",
				"101111101111",
				"101111101110",
				"101011011110",
				"011110011010",
				"100010101011",
				"100111011101",
				"101011101110",
				"101111101111",
				"100111001101",
				"100110111100",
				"100111001101",
				"101011011110",
				"101111101111",
				"100110111101",
				"011110101011",
				"101011011111",
				"101011101111",
				"101011111111",
				"100111101111",
				"100111011110",
				"101111101111",
				"110011101111",
				"011010001001",
				"010101111000",
				"100111001101",
				"100111101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101111101111",
				"011110011011",
				"011010001001",
				"101011011110",
				"101111101111",
				"110011111111",
				"110011101111",
				"100110111101",
				"011110011011",
				"011110101100",
				"011111011110",
				"100011101110",
				"100011101111",
				"101011101111",
				"110011011111",
				"101010111100",
				"011110011011",
				"100011001101",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"011111101111",
				"011111111111",
				"100011101111",
				"100111101111",
				"100111011111",
				"100011011111",
				"011111011111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011011110",
				"011110111100",
				"101011001101",
				"110011001110",
				"100010001001",
				"011001100111",
				"100110101100",
				"100110111101",
				"100011001110",
				"011111011110",
				"011011011111",
				"011011101111",
				"011111011111",
				"011111011110",
				"100011001110",
				"100011001110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011110",
				"010010101011",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"011110111100",
				"011010011011",
				"011010011010",
				"100110101100",
				"101111001101",
				"110011001110",
				"101111001110",
				"101010111101",
				"100110111101",
				"011110101100",
				"011110111101",
				"100011001110",
				"010110101100",
				"011010111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111010",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"011110101010",
				"100010101011",
				"010101100110",
				"010101000110",
				"100010001001",
				"100010011010",
				"011010101010",
				"010110101010",
				"011010101011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011110111011",
				"011110111011",
				"011010101011",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110101010",
				"011010111011",
				"010110101010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110101001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010011001",
				"010101111000",
				"001101010101",
				"001000110100",
				"001100110100",
				"010001010110",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001001",
				"010101110111",
				"010001100110",
				"011001111000",
				"011110011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110000111",
				"010101110111",
				"010101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010011001",
				"011010011001",
				"010110001001",
				"010001111000",
				"001101110111",
				"001101110111",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010001110111",
				"001101100111",
				"001101100111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"110011001011",
				"101111001011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110111011110",
				"110111011110",
				"110111011110",
				"110111011101",
				"110111001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101011001110",
				"101011001110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111101110",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011110",
				"101111011110",
				"101011011101",
				"101011011101",
				"101011011110",
				"101111101110",
				"101111011110",
				"101111001101",
				"101011001101",
				"101111101110",
				"110011101111",
				"110011101110",
				"110011011110",
				"101111001101",
				"100110111100",
				"101011001101",
				"101111101110",
				"110011101111",
				"101111101110",
				"101011011101",
				"100010101011",
				"100110111100",
				"101011011110",
				"101011101110",
				"101111011110",
				"100010101011",
				"011110011011",
				"100110111101",
				"101111101111",
				"101111101111",
				"100010111100",
				"011110101011",
				"101111011111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111011110",
				"011110001001",
				"011010001001",
				"100111011110",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111111111",
				"100011111111",
				"101111101111",
				"100110111100",
				"010101111000",
				"100110101100",
				"110011011111",
				"101111001110",
				"100010101100",
				"100010011011",
				"100010101100",
				"100111001110",
				"100011011110",
				"011111101110",
				"100011101110",
				"100111101111",
				"110011111111",
				"101011001110",
				"011010001010",
				"100011001101",
				"100011101111",
				"011011011110",
				"100011101111",
				"011111101111",
				"011111111111",
				"011111111111",
				"100011101111",
				"100111101111",
				"100111011111",
				"100111101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111001101",
				"100011001101",
				"101111011110",
				"110011011110",
				"100110011011",
				"011110001001",
				"100010011010",
				"100010111100",
				"100010111101",
				"011111011110",
				"011111011111",
				"011011101111",
				"011011011111",
				"011111011111",
				"011111001110",
				"011111001110",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011111001100",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001100",
				"011111001101",
				"011111001101",
				"100011011101",
				"100011011110",
				"011010101011",
				"011110111100",
				"100011001101",
				"100111011110",
				"100111011110",
				"101011011111",
				"101011101111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100010101101",
				"011110101100",
				"011010011011",
				"010110011011",
				"011010111100",
				"011111001101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011101111",
				"101011101111",
				"011110111101",
				"011010011011",
				"011110101100",
				"100010111101",
				"011110111100",
				"011010101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010111001011",
				"010111001011",
				"011010111011",
				"011110111011",
				"011110101011",
				"011010111011",
				"010110111011",
				"010110111010",
				"011110111011",
				"011110101010",
				"011110001000",
				"011001100111",
				"011001111000",
				"011110011010",
				"011110111011",
				"010110111011",
				"010110111011",
				"011010111100",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011110111011",
				"011010101010",
				"010110011001",
				"011010101010",
				"011010111011",
				"011110111011",
				"010110101010",
				"010010001000",
				"010110101010",
				"010110101010",
				"010110011001",
				"010010011001",
				"010110101010",
				"011010111010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011110111011",
				"011110111011",
				"010110011001",
				"010010001000",
				"001101110111",
				"001101100111",
				"010001100111",
				"010001100111",
				"010101100111",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010001111000",
				"010110001000",
				"011010001001",
				"011110001001",
				"011110001000",
				"011010001000",
				"011010001001",
				"011010011010",
				"010110001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010010000111",
				"010001110111",
				"010010001000",
				"010010000111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010011001",
				"011010001001",
				"010110001000",
				"010001110111",
				"001101110111",
				"001101100110",
				"001101100111",
				"010001110111",
				"010110001000",
				"010110001000",
				"010110001000",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001001",
				"010001111000",
				"010001110111",
				"010001111000",
				"010101111000",
				"010001111000",
				"010001111000",
				"010110001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011010",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011101111",
				"110011101111",
				"110011011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011001101",
				"100111001101",
				"100111001100",
				"101011011110",
				"101011011110",
				"101011101110",
				"101011101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101111101110",
				"110011101111",
				"101111101110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101011001101",
				"101011011101",
				"101111101110",
				"101111101110",
				"101111011110",
				"101111001110",
				"101011011101",
				"101111101110",
				"101111011110",
				"101111011110",
				"110011011110",
				"101111001101",
				"101011001101",
				"101011011101",
				"101111101110",
				"110011101111",
				"110011101111",
				"101111001101",
				"100010101011",
				"100111001100",
				"101011101110",
				"101011101111",
				"101111011110",
				"011110001001",
				"011110001010",
				"100111001101",
				"101111101111",
				"101111101111",
				"011110101011",
				"011110101011",
				"101111101111",
				"101011011110",
				"101011101110",
				"101111101111",
				"101111101111",
				"101111011110",
				"100010011010",
				"011001111000",
				"011110011011",
				"101011011110",
				"100111101111",
				"100111101111",
				"100011101111",
				"011111111111",
				"100011111111",
				"100011111111",
				"101011101111",
				"101011001101",
				"010101101000",
				"011001101000",
				"100110011011",
				"100010011011",
				"011110011011",
				"100110111101",
				"100111011110",
				"100111011111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111011110",
				"101011101111",
				"101111101111",
				"100010101011",
				"011110111100",
				"011111001101",
				"011111011110",
				"100011101111",
				"100011101111",
				"011111111111",
				"011111101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100011101111",
				"100011101110",
				"100111101111",
				"100111101111",
				"101011011111",
				"110011101111",
				"101010111101",
				"011110001001",
				"011110001001",
				"100010011011",
				"100111001110",
				"100011001110",
				"011111011110",
				"011011101111",
				"011011101111",
				"011011011111",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100011001101",
				"011110111100",
				"011110111100",
				"101011101111",
				"011010101011",
				"011110101011",
				"100110111101",
				"101011001110",
				"101011001110",
				"100110111101",
				"100010111100",
				"100010101100",
				"011110101011",
				"011010011011",
				"011110011100",
				"011110101100",
				"011110101100",
				"011110111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011011001101",
				"011111011110",
				"100111101111",
				"100111011110",
				"100010111101",
				"011110101100",
				"011110101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010010111011",
				"010010111011",
				"010110111011",
				"011010101011",
				"011010101011",
				"011010111011",
				"010110111011",
				"010110111010",
				"010110101010",
				"011110101010",
				"100110101011",
				"100001111000",
				"011001100111",
				"011110011010",
				"011010111011",
				"010010111010",
				"010110111011",
				"010110111100",
				"010110111011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010101001",
				"010010101001",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010111011",
				"011010101010",
				"010110101010",
				"010010001001",
				"010110011001",
				"011010101010",
				"011010101010",
				"010110101001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011110111011",
				"011110111011",
				"011010101010",
				"010110011001",
				"010010001000",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001111000",
				"010110001001",
				"011010011001",
				"011110011010",
				"100010011010",
				"100010101011",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"011010101010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110011001",
				"010110001001",
				"010101110111",
				"010101111000",
				"011110001001",
				"011110001001",
				"011001111000",
				"010101111000",
				"011010001001",
				"010110001001",
				"010001111000",
				"010110011001",
				"010110011010",
				"010010001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010110001000",
				"010001110111",
				"010101111000",
				"010001110111",
				"010101111000",
				"010110001000",
				"010001110111",
				"001101100111",
				"001101100111",
				"001101110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"010110001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001111000",
				"010110001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"000100010010",
				"001000100010",
				"001100110100",
				"010001000100",
				"010101010101",
				"010101100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110111011101",
				"110111011101",
				"110111011101",
				"110111001101",
				"110111001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111101110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011001101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101111011110",
				"101111101110",
				"101111101111",
				"101111101110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111101110",
				"101111101110",
				"110011011110",
				"101111011110",
				"101011001101",
				"101111011110",
				"101111001101",
				"101111001101",
				"110011011110",
				"101111011101",
				"101011011101",
				"101111011110",
				"110011101111",
				"110011101111",
				"110011011110",
				"101010111100",
				"100110101011",
				"100111001101",
				"101011101110",
				"101111101111",
				"101011001101",
				"011001111001",
				"011110001010",
				"101011001110",
				"101111111111",
				"101011101111",
				"011010011011",
				"100010111100",
				"101111101111",
				"101111101111",
				"101011101111",
				"101111101111",
				"101111101110",
				"101011001101",
				"011101111001",
				"011101111000",
				"100110111100",
				"101011011110",
				"101011101111",
				"100111111111",
				"100011111111",
				"100011111111",
				"011111111111",
				"100111111111",
				"100111101110",
				"101111011110",
				"100010001010",
				"010101010111",
				"011101111001",
				"100010011010",
				"101011001110",
				"100111001110",
				"100111011110",
				"100111101111",
				"100111101111",
				"100011101111",
				"011111101110",
				"011111011110",
				"100011011110",
				"101111111111",
				"101011011110",
				"011010011011",
				"011111001101",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"100111101111",
				"100111011111",
				"100111101111",
				"101011101111",
				"100111011110",
				"101111101111",
				"101011011110",
				"100110111100",
				"011110001010",
				"011110001001",
				"100110101100",
				"100110111100",
				"100111001110",
				"011111001110",
				"011111011111",
				"011111101111",
				"011011101111",
				"011011011111",
				"011111011111",
				"100011011111",
				"100011001110",
				"011111001101",
				"011011011101",
				"011011011101",
				"011011011101",
				"011111001101",
				"011111001100",
				"100010111100",
				"011110111101",
				"100011001110",
				"100011001101",
				"100011001101",
				"011111001101",
				"011110101011",
				"101011011110",
				"011110011011",
				"011001111001",
				"011101111001",
				"011101111001",
				"011101111010",
				"011110001011",
				"100010011100",
				"100010101100",
				"011110101100",
				"011110101100",
				"011110111101",
				"011111011110",
				"011111011110",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001110",
				"100011001110",
				"011111001110",
				"011111001110",
				"011011001101",
				"011111011110",
				"100111101111",
				"100011011110",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"011010101010",
				"100110111011",
				"101010101011",
				"011001100111",
				"011001101000",
				"011110101010",
				"010110101010",
				"010010101010",
				"010110111100",
				"010110111100",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101001",
				"010010101001",
				"010010101001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011010",
				"011010101010",
				"011110111011",
				"011010101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"011010011010",
				"011010011001",
				"011110101010",
				"100010111011",
				"011110111011",
				"011110101010",
				"011010011010",
				"010010001000",
				"001101110111",
				"001001100110",
				"001101110111",
				"001101110111",
				"001110001000",
				"010010001000",
				"010110011001",
				"011010011010",
				"011010011001",
				"011010001001",
				"011110011010",
				"100010101011",
				"011110101010",
				"011010011010",
				"010110011001",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110001001",
				"010001110111",
				"010101110111",
				"011110001001",
				"011110001001",
				"011001111000",
				"010101100111",
				"011010001001",
				"011010001001",
				"010101111000",
				"010110001001",
				"010110011001",
				"010010001001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010001000",
				"010010000111",
				"010010000111",
				"010010000111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"001101100110",
				"010001100111",
				"010001110111",
				"010101111000",
				"010101110111",
				"010001100111",
				"010101110111",
				"010101110111",
				"010101111000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010010001000",
				"001101110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101100111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010110001000",
				"010110001000",
				"010101111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"000100100010",
				"001000110011",
				"001100110100",
				"010001000101",
				"010101010101",
				"010101010110",
				"011001100110",
				"011001100111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011010",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101001",
				"101110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110111001101",
				"110111001101",
				"110111001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111101110",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111011111",
				"110011011111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011101110",
				"101111101111",
				"101111101110",
				"101111101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"100110111101",
				"101010111101",
				"101011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"101111011110",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111011110",
				"110011101110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"110011011110",
				"101111011110",
				"101011011101",
				"101111101110",
				"110011101111",
				"110011011110",
				"110011001110",
				"101010101100",
				"100110111100",
				"101011011110",
				"101011101110",
				"101111101111",
				"101011001101",
				"011010001001",
				"100010011011",
				"101111011110",
				"101111101111",
				"101011101111",
				"011010011010",
				"011110101011",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101111011110",
				"011110001001",
				"100010001010",
				"101011001101",
				"101011011110",
				"101011101111",
				"101011101111",
				"100111111111",
				"100011111111",
				"100011101111",
				"100111111111",
				"100111011110",
				"110011101111",
				"101110111100",
				"011001010111",
				"011101111001",
				"100110111100",
				"100011001101",
				"100011011111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101110",
				"101011101111",
				"101011101111",
				"011010101011",
				"011110111101",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011011110",
				"100010101011",
				"011001111001",
				"011110001010",
				"100110101011",
				"100110101100",
				"101010111101",
				"100010111100",
				"100011001110",
				"011111001110",
				"011111011111",
				"011011101111",
				"011111101111",
				"011111011111",
				"011111011110",
				"100011011110",
				"100011001110",
				"011111011101",
				"011111011101",
				"011011101101",
				"011111101110",
				"011111011101",
				"100011001101",
				"100010111101",
				"100010111101",
				"011110111101",
				"011110111101",
				"100011011110",
				"011111001100",
				"011010111011",
				"100111011110",
				"100110111100",
				"100010011010",
				"011101111001",
				"100001111001",
				"101010011100",
				"100110101101",
				"100010101100",
				"100010101101",
				"011110111101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011110111101",
				"011111001110",
				"100011011111",
				"011011001101",
				"011011001101",
				"011111011110",
				"011111011110",
				"011111001101",
				"011010111011",
				"011010111011",
				"011010111100",
				"011110111100",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011011001011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"100010111011",
				"011001111000",
				"011001100111",
				"010101010110",
				"011001111000",
				"011110011010",
				"011010101011",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101010",
				"010110011001",
				"010110001000",
				"011010011001",
				"100010101011",
				"100010101011",
				"011110011001",
				"010101110111",
				"001101100111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110011001",
				"010010011001",
				"010110011001",
				"010110011010",
				"011010011001",
				"010110001001",
				"010110001001",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110001000",
				"011010001000",
				"011110001000",
				"011001111000",
				"011001100111",
				"010101100111",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101110111",
				"010101111000",
				"010101111000",
				"010101111000",
				"011010001001",
				"011010001000",
				"011010001001",
				"010110001001",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010010001000",
				"010001110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010101111000",
				"011010001001",
				"011010001000",
				"010101110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000110011",
				"001100110100",
				"010001000100",
				"010001010101",
				"010101010110",
				"011001100110",
				"011001100111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110111011110",
				"110011011110",
				"110011011110",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011011111",
				"110011011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011101111",
				"101111101111",
				"101111011111",
				"110011101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011001110",
				"101010111101",
				"101010111101",
				"101111011110",
				"101111011111",
				"101111011110",
				"101111011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"101011001101",
				"101010111100",
				"101111001101",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101011001101",
				"101011001101",
				"101111001101",
				"110011011110",
				"110111101111",
				"101111011101",
				"101011011101",
				"101111101110",
				"110011101110",
				"110011001110",
				"110111001110",
				"101110111100",
				"101011001101",
				"101011011110",
				"101011101110",
				"101111101111",
				"101011001101",
				"011010001001",
				"100110111100",
				"101111011110",
				"101011101111",
				"101011101111",
				"011010011011",
				"011110101011",
				"101011101111",
				"101111101111",
				"101011101111",
				"101011011110",
				"110011101111",
				"110111101111",
				"100110011010",
				"100010011010",
				"101011011110",
				"101011011110",
				"101111101111",
				"101011101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011101110",
				"110011101111",
				"110011001110",
				"011001101000",
				"011110001001",
				"100111001101",
				"011111001101",
				"011111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100011011110",
				"100011101111",
				"100011101111",
				"101011111111",
				"011110111101",
				"011010101100",
				"100111011110",
				"100011101111",
				"100011101110",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"100111001101",
				"100010101100",
				"101011001101",
				"110011001110",
				"110011001110",
				"101010111101",
				"100110101100",
				"100110111100",
				"100111001101",
				"100010111101",
				"011111001110",
				"011111011111",
				"011011101111",
				"011011101111",
				"011111011111",
				"100011011110",
				"100011001110",
				"100011001101",
				"011111011101",
				"011111011101",
				"011011101101",
				"011111101110",
				"011111101110",
				"100011011110",
				"100011001110",
				"100011011111",
				"011010111101",
				"011011001101",
				"011111011110",
				"010111001100",
				"100011101110",
				"011111001100",
				"100111001100",
				"100010101010",
				"011001101000",
				"011101111001",
				"101010111101",
				"101011001101",
				"100010111101",
				"011110111101",
				"011111001101",
				"100011001110",
				"100011011110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011111011101",
				"011111001101",
				"100011011110",
				"011110111100",
				"011110111011",
				"011010111100",
				"011010111100",
				"011111001101",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011011001100",
				"011111001100",
				"011111001100",
				"011111001011",
				"011111001011",
				"011110111011",
				"011110111011",
				"011110111011",
				"011110101011",
				"011110111100",
				"011110101011",
				"011110101011",
				"011110011010",
				"011010001000",
				"001000110100",
				"010001000101",
				"100001111001",
				"100010001010",
				"100010011011",
				"011110111100",
				"010110111011",
				"010110111100",
				"010110111100",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010101011",
				"010110101010",
				"011010101010",
				"011010111010",
				"010110111010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011110101011",
				"011010011010",
				"010001100111",
				"001001000100",
				"001000110100",
				"010001010101",
				"010101100110",
				"010101100111",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"011010011010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010011010",
				"011010011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011010001000",
				"010101100111",
				"011001100111",
				"011101111000",
				"010101111000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011000",
				"010110011000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101110111",
				"010101110111",
				"010101110111",
				"011001111000",
				"011110001001",
				"011001111000",
				"010101111000",
				"011010011001",
				"010001111000",
				"010010001000",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"001101110111",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"001101110111",
				"001101100110",
				"001101100110",
				"010001110111",
				"010101111000",
				"010101110111",
				"010001100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011000",
				"101010011000",
				"101010011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110010111100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110111011101",
				"110111011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111101111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011011111",
				"110011101111",
				"110011011111",
				"110011011110",
				"101111011110",
				"101111011101",
				"110011011110",
				"110011101110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111011111",
				"101011001110",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111101111",
				"101111101111",
				"101111011110",
				"101010111101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"110011101110",
				"110011101111",
				"110011011110",
				"110011011110",
				"101011001101",
				"101011001100",
				"101111001101",
				"110011101110",
				"110111101111",
				"101011001101",
				"101011011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"110111011110",
				"110011001101",
				"101111011101",
				"101011011110",
				"101111101110",
				"110011101111",
				"101011001100",
				"011110011010",
				"101011001101",
				"101111101111",
				"101011011110",
				"101111101111",
				"011110101011",
				"100110111100",
				"101111101111",
				"101011011110",
				"100111001101",
				"100111001101",
				"110011101111",
				"110111101111",
				"100110101011",
				"011110011010",
				"100111011101",
				"100111101110",
				"101111101111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"101011101111",
				"110011101111",
				"110111011110",
				"011001101000",
				"011010001010",
				"100011001101",
				"100011101110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"101011111111",
				"100111011110",
				"010110001010",
				"100111001110",
				"101011111111",
				"100011011110",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111111111",
				"101011101111",
				"100011001101",
				"011110101011",
				"011010011010",
				"100010111100",
				"101011001110",
				"110011011111",
				"110111101111",
				"110111101111",
				"101111001110",
				"100110111100",
				"100010111101",
				"100011001110",
				"100011001111",
				"011111011111",
				"011011011110",
				"011011011110",
				"011111011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111101110",
				"011111101110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011011111",
				"011111101111",
				"011011001101",
				"011011011101",
				"011011011100",
				"011111001100",
				"011111001100",
				"100111001101",
				"011010001001",
				"011110001010",
				"100110111101",
				"100110111101",
				"100010111101",
				"100011011110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011011001110",
				"011011001110",
				"011011001101",
				"011011001110",
				"011111011110",
				"010111001101",
				"011011001100",
				"011111001101",
				"011110111100",
				"100011001101",
				"100011001101",
				"011110111100",
				"011010111011",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110001000",
				"001101010110",
				"010001010110",
				"011001100111",
				"011101111001",
				"100010011010",
				"100010101011",
				"011110111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010111010",
				"011010111010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"010110101010",
				"010110011001",
				"011010011001",
				"100010101011",
				"011110011010",
				"010001100110",
				"001101000100",
				"010101010110",
				"011110001001",
				"100010011010",
				"011010011001",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110101010",
				"010110011010",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"011010001000",
				"011001111000",
				"011001111000",
				"011001111000",
				"010110001000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010010011001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001110000111",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010101111000",
				"011010001000",
				"011001111000",
				"011001111000",
				"011010001001",
				"011001111000",
				"010101111000",
				"010110011001",
				"010001111000",
				"010010001000",
				"010110011001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"001101110111",
				"001101100111",
				"001101100111",
				"010001100111",
				"010001100111",
				"010101110111",
				"010101111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011110000111",
				"100010001000",
				"100010001000",
				"100010001001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010011000",
				"101010011000",
				"101010011000",
				"101010011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011011111",
				"101111011110",
				"101111011111",
				"101111101111",
				"101111101111",
				"101111011110",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101110",
				"101111011110",
				"101011001101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011101111",
				"110011011110",
				"101111011110",
				"101011001101",
				"101111001101",
				"101111011110",
				"110011011110",
				"110011101111",
				"101111011110",
				"101111011101",
				"101011001101",
				"101111001101",
				"101111001101",
				"110011011110",
				"110011011110",
				"101111001101",
				"101111011101",
				"110011101110",
				"110111101111",
				"100110111011",
				"100010101011",
				"101011011110",
				"101011101111",
				"101111101111",
				"101111011111",
				"100010011010",
				"101010101100",
				"101111011110",
				"100110111100",
				"100111011101",
				"100111011110",
				"101111101111",
				"110011101111",
				"100010011010",
				"011110011010",
				"100111101110",
				"100111111111",
				"100111111111",
				"100111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011011101",
				"101111101111",
				"110111111111",
				"101010101100",
				"011001111001",
				"011010011011",
				"100011011110",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111111111",
				"011010011011",
				"100111001101",
				"110111111111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011011111",
				"100110111101",
				"011110101011",
				"011010101011",
				"011110111101",
				"100011001110",
				"100111011111",
				"100111011111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"100111001101",
				"011010101011",
				"100111001111",
				"011110111110",
				"100011101111",
				"011111011111",
				"011011001110",
				"011111011110",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100111011111",
				"100011001110",
				"011111001110",
				"011111011110",
				"011111101110",
				"011011011101",
				"011111011101",
				"100011011101",
				"100111011101",
				"010110001001",
				"011110011010",
				"100110101101",
				"100010111101",
				"100011001110",
				"011010111110",
				"011111011111",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"100011011101",
				"011010111011",
				"010110101010",
				"011111001101",
				"011111001101",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001100",
				"100011001100",
				"100010111100",
				"100011001100",
				"011110111100",
				"011110111100",
				"011010101011",
				"010010001001",
				"010001111000",
				"010110001001",
				"011110101011",
				"100111001101",
				"101011011110",
				"101011001101",
				"100010111100",
				"011110011010",
				"011010001001",
				"011110011011",
				"011110111100",
				"011110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110111010",
				"010110011001",
				"011010011001",
				"100010101010",
				"011110001000",
				"010101010110",
				"010101110111",
				"011010001000",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011010011001",
				"011010011001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010001111000",
				"010001110111",
				"010101111000",
				"011010001001",
				"011010001001",
				"011010011001",
				"011110011010",
				"011010101010",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010001111000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"010101111000",
				"010001110111",
				"010101110111",
				"010101110111",
				"011001111000",
				"011110001001",
				"011010001000",
				"010001110111",
				"010010001000",
				"010010001000",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010001111000",
				"010010001000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010110",
				"010101100110",
				"011001110111",
				"011101110111",
				"011101111000",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011000",
				"101010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011111",
				"110011011110",
				"110011011110",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"101111011110",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"101010111100",
				"101011001101",
				"101111011110",
				"110011101110",
				"110011101111",
				"101111011110",
				"101111001110",
				"101010111100",
				"101111001101",
				"101111011101",
				"110011011110",
				"110011011110",
				"101111011101",
				"110011101110",
				"110011101110",
				"110011101110",
				"101010111011",
				"100110101011",
				"101011011110",
				"101011101111",
				"101011101111",
				"101111101111",
				"011101111001",
				"100001111001",
				"100110101011",
				"100010111011",
				"100111011101",
				"100111101110",
				"101111111111",
				"110011111111",
				"100010101011",
				"011010001010",
				"011111001101",
				"100011101110",
				"100011111111",
				"101011111111",
				"101111101111",
				"101111011111",
				"101111011110",
				"110011101111",
				"110011101110",
				"100110111100",
				"011101111001",
				"011110001010",
				"100010111101",
				"100011011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011110",
				"101011101111",
				"011010011010",
				"011010001010",
				"101010111101",
				"101010111101",
				"101110111101",
				"101010101100",
				"100010011011",
				"011110011011",
				"011110101100",
				"100011001110",
				"100111011111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011011110",
				"011110111100",
				"100011001110",
				"011111001111",
				"100011011111",
				"100011101111",
				"011111011110",
				"100011101111",
				"100011011111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011111",
				"100111011111",
				"100011011111",
				"100011011110",
				"011111011110",
				"100011011111",
				"100111001111",
				"100111011111",
				"100111011111",
				"100011011110",
				"011111011101",
				"011111011101",
				"100011011101",
				"100111011101",
				"100111001101",
				"011010001001",
				"011010001010",
				"100010101100",
				"100010111110",
				"100011001111",
				"011111001111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011111001101",
				"011010111100",
				"100011001101",
				"011111001100",
				"010110011010",
				"011110111100",
				"100111011110",
				"100011001101",
				"100011001101",
				"100111001110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001100",
				"011110101011",
				"011010101011",
				"010110011001",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111011",
				"011111001100",
				"100011001101",
				"011110111100",
				"100011001101",
				"100011001101",
				"100111011110",
				"100011001101",
				"011010101011",
				"011010011010",
				"011010101011",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010010101010",
				"010010111010",
				"011010111010",
				"010110011001",
				"100010011010",
				"100010011001",
				"011001110111",
				"010101100111",
				"010110001000",
				"010110101001",
				"010010011010",
				"010010011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"010110011001",
				"011010011001",
				"011110101010",
				"011110011010",
				"011110101010",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110001001",
				"010001111000",
				"001101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"011010011010",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010011001",
				"010110011001",
				"010010001000",
				"001110001000",
				"010010001000",
				"010110001001",
				"011010011001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010101111000",
				"011010001000",
				"011010001001",
				"011010001000",
				"010001110111",
				"010110001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101111000",
				"001101111000",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001110111",
				"010101111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001000",
				"010110001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110011",
				"001101000100",
				"010001010101",
				"010101010110",
				"011001100110",
				"011001100111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011000",
				"101010011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110111011110",
				"110111011110",
				"110111011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011111",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"101011001101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111001110",
				"101010111100",
				"101011001101",
				"110011011110",
				"110011101110",
				"110011011110",
				"101111011101",
				"110011101110",
				"110011101110",
				"101111011101",
				"101010111100",
				"101010111100",
				"101111101111",
				"101111101111",
				"101011011110",
				"110011101111",
				"011101111001",
				"011001100111",
				"011110001001",
				"100010111011",
				"100011011101",
				"100111101110",
				"101111111111",
				"110011101111",
				"100010011010",
				"011110001001",
				"100111011110",
				"100111101111",
				"100111111111",
				"100111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111101110",
				"100111001100",
				"011110001001",
				"011001111000",
				"100010011011",
				"100111001110",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011001101",
				"101011101111",
				"100010111100",
				"010101111000",
				"100010001010",
				"100110011011",
				"011110001010",
				"100010011011",
				"100010101100",
				"100110111101",
				"100111011110",
				"100111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"011110111101",
				"011111001110",
				"011111011111",
				"100011101111",
				"011111011111",
				"100011111111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100111101110",
				"101011101111",
				"101011011101",
				"100110111100",
				"011010001001",
				"011110001001",
				"100010011011",
				"100010111101",
				"100011001110",
				"011111001110",
				"011011011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001101",
				"011010111100",
				"011111001101",
				"100011001101",
				"011110111011",
				"011110101011",
				"100010101100",
				"100110111101",
				"100110111101",
				"100110111101",
				"100010101100",
				"011010011011",
				"011010011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110101010",
				"011010111100",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011110111100",
				"011111001100",
				"100011011101",
				"100011011101",
				"011111001101",
				"011010111011",
				"010110011010",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010011001",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110111010",
				"010110101010",
				"010110011000",
				"100010011010",
				"100110011010",
				"011101111000",
				"010101110111",
				"010110001000",
				"011010101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"011110101011",
				"011110101011",
				"011010011010",
				"011110101010",
				"011110011010",
				"010110001001",
				"010001111000",
				"001101111000",
				"001101111000",
				"010001111001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001001",
				"010010001000",
				"010010001001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010001110111",
				"010110001000",
				"010110001000",
				"011010001001",
				"011010001000",
				"010101110111",
				"010001100111",
				"010101110111",
				"010110001000",
				"001101110111",
				"010001110111",
				"010110001000",
				"010110011001",
				"010010001000",
				"001101110111",
				"001101111000",
				"010010001000",
				"001101111000",
				"001101111000",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001110111",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001010101",
				"010101010110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100001111000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110111011110",
				"110111011110",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"101010111101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111001110",
				"101010111100",
				"101111001101",
				"110011011110",
				"110011101110",
				"101111011101",
				"101111001101",
				"110011011110",
				"101111011101",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111101111",
				"101111101111",
				"101011011110",
				"110011101111",
				"100110011010",
				"011001100111",
				"011110001001",
				"101011011101",
				"100111101110",
				"100111101110",
				"101011101111",
				"101111101111",
				"100010011010",
				"100010001010",
				"101011011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"101111101111",
				"110011101111",
				"101111101110",
				"101011011101",
				"100110111100",
				"100010011010",
				"100010001010",
				"100110101100",
				"100111011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100111101111",
				"100111011110",
				"101011101111",
				"101111011110",
				"011110001010",
				"011101111001",
				"100110011011",
				"100110101011",
				"100110111101",
				"101011011110",
				"101011011111",
				"100111011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"011111011111",
				"011111011110",
				"100011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111111111",
				"100011001110",
				"011010111101",
				"011111011110",
				"011111011110",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101110",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111011110",
				"101011011110",
				"101011001100",
				"100010011010",
				"011001100111",
				"011001100111",
				"100110011011",
				"100110101100",
				"100010111101",
				"100011001110",
				"011011001110",
				"011011011111",
				"011011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"010111001100",
				"011011001101",
				"011010111100",
				"011111001100",
				"100111011101",
				"100010101011",
				"011010001001",
				"100010011011",
				"011110001010",
				"011110011010",
				"011010001010",
				"011010001010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011110111100",
				"011111001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011010111100",
				"010110011010",
				"011010101011",
				"011010101011",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010111011",
				"011110111011",
				"011110101011",
				"011110101010",
				"011110101011",
				"011010101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011110101010",
				"100110101011",
				"100010001001",
				"010101010110",
				"010101100110",
				"010110001000",
				"011010101010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011000",
				"010010011000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"010010001000",
				"001101100111",
				"001101100111",
				"010101111000",
				"011010001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010001111000",
				"010001111000",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010110001001",
				"001101111000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"011010011001",
				"010110001000",
				"010101111000",
				"010101111000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"001101110111",
				"001101110111",
				"010010001000",
				"010110001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"001101110111",
				"001101110111",
				"001101110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"010001110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000010001",
				"000100010010",
				"001000100010",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100001111000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"110011001100",
				"110011001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110111011101",
				"110011011101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011101",
				"101011001101",
				"101111011101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"101010111100",
				"101111001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101011001101",
				"101010111100",
				"101111011110",
				"110011101110",
				"110011011110",
				"101111011110",
				"101111001101",
				"101011001101",
				"101011001100",
				"101111001101",
				"110011011110",
				"101111001110",
				"101111011110",
				"101111101111",
				"101011011110",
				"110011011110",
				"100110011010",
				"011001100111",
				"100010011010",
				"101111101110",
				"100111101110",
				"100111101110",
				"101011101111",
				"110011101111",
				"100110101011",
				"100010011010",
				"101011001110",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111101111",
				"101111011110",
				"100010111100",
				"101011011110",
				"101111101110",
				"101010111100",
				"100110011011",
				"100110101100",
				"101011011111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100111101111",
				"101011101110",
				"101111101111",
				"100110111100",
				"011001111000",
				"100010011011",
				"101011001101",
				"101011011110",
				"100111011110",
				"100111011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111011111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"011110111101",
				"011111001110",
				"100011101111",
				"100011101111",
				"011111101110",
				"100011111111",
				"011111101110",
				"100011111111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011110",
				"100011101110",
				"100111101111",
				"101011101111",
				"100111001101",
				"011010001001",
				"010001010110",
				"010101010110",
				"011001100111",
				"100010001001",
				"101010111100",
				"100110101100",
				"100010111100",
				"100011011110",
				"011111011110",
				"011111101111",
				"011011011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011111001100",
				"011111001100",
				"100010111100",
				"100110111100",
				"100010011010",
				"010101100111",
				"011110001010",
				"011110011011",
				"011110101011",
				"100010101100",
				"100010111101",
				"100010111101",
				"100010111101",
				"100011001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001100",
				"011010111100",
				"010110111011",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"100011011101",
				"100011011101",
				"011010011010",
				"010110011010",
				"010110101010",
				"011010111011",
				"011010111100",
				"011010111100",
				"010110111100",
				"010111001100",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111010",
				"011010111011",
				"011010001001",
				"010101100111",
				"010001000101",
				"010101000110",
				"011101111000",
				"011110011010",
				"011110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110001001",
				"010110011001",
				"010001100111",
				"001001000101",
				"010001100110",
				"011110011010",
				"011010001001",
				"011010011001",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010110101011",
				"010110011010",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010010001001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110001000",
				"010001100111",
				"001101100111",
				"010001110111",
				"010110001000",
				"010110001000",
				"011010011001",
				"010110011001",
				"011010011001",
				"010110001001",
				"010001111000",
				"001101110111",
				"010001111000",
				"010110001001",
				"010010001001",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010101111000",
				"010101111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100001111000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011001101",
				"110011011110",
				"110011011110",
				"101111011110",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111001101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011110",
				"101111011110",
				"110011011110",
				"101111001101",
				"101011001100",
				"101111011101",
				"101111011110",
				"101011011101",
				"101111011110",
				"101111011110",
				"101010111100",
				"100110111100",
				"101111011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111001101",
				"100110111100",
				"101011001100",
				"101111011110",
				"110011011111",
				"101111011110",
				"101111011110",
				"101111101110",
				"101111011110",
				"110011011110",
				"100010001001",
				"011001100111",
				"100010101011",
				"101111101110",
				"100111101110",
				"100011101110",
				"101011101111",
				"101111101111",
				"101010101011",
				"100110011010",
				"101111001110",
				"110011101111",
				"110011111111",
				"101111101111",
				"101011011110",
				"100010111100",
				"100011001100",
				"101011011110",
				"110011111111",
				"101111011110",
				"100110011011",
				"100110101101",
				"101011011111",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100011111111",
				"100011101111",
				"100111101111",
				"100111011110",
				"101111101111",
				"101111011101",
				"011001111000",
				"100010011011",
				"100111001101",
				"100111011110",
				"100111011110",
				"100111011111",
				"100111101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011011111",
				"100011011110",
				"101111111111",
				"100011001110",
				"011111001101",
				"100111101111",
				"100011011110",
				"100111101111",
				"100111111111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"100111101111",
				"011010111100",
				"010010001001",
				"011010011010",
				"100010101011",
				"100110101011",
				"100110011010",
				"100010001001",
				"100010001010",
				"101010101100",
				"100010111100",
				"100011001101",
				"100011011110",
				"011111011110",
				"011111101111",
				"011011011111",
				"011011011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"010110111100",
				"011111001101",
				"100011001101",
				"011110101011",
				"100110111100",
				"100110111100",
				"011010001000",
				"100010101011",
				"100010101100",
				"100010101100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001100",
				"011111001100",
				"011010111011",
				"011110111100",
				"011010101011",
				"010110011010",
				"010110101010",
				"011010111100",
				"011011001100",
				"010111001100",
				"010110111100",
				"010111001100",
				"010111001100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101010",
				"011010111011",
				"011010111011",
				"010110111010",
				"010110101010",
				"010110011001",
				"010001100111",
				"001101000110",
				"010001000101",
				"011001010111",
				"100010001001",
				"011110001001",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101001",
				"010110101001",
				"011010101010",
				"011010011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"011010011001",
				"011010011001",
				"010101111000",
				"011001111000",
				"011110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010010011001",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010010011001",
				"010010001001",
				"010010011001",
				"010110011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110011001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010110001001",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"010110011010",
				"010010001000",
				"001101110111",
				"001101100111",
				"001101100111",
				"010001111000",
				"010110001000",
				"010001110111",
				"010001110111",
				"010010001000",
				"010110001001",
				"011010011001",
				"011010011010",
				"010110001001",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100011",
				"001100110011",
				"010001000100",
				"010101000100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101111000",
				"100010001000",
				"100010001000",
				"100010011001",
				"100010011001",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"110011001100",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011101",
				"101111011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"101111011101",
				"110011011110",
				"101111011101",
				"101011001101",
				"101111001101",
				"101111011110",
				"101011001101",
				"101111011110",
				"101011001101",
				"100110111100",
				"100110111100",
				"101111001101",
				"110011011110",
				"101111011110",
				"110011011110",
				"101111001101",
				"100110111100",
				"101011001101",
				"110011011110",
				"110011011110",
				"101111011110",
				"101111011101",
				"101111011110",
				"110011101110",
				"110011011101",
				"100010001000",
				"011101111000",
				"101010111100",
				"101111101110",
				"100111111111",
				"100011101110",
				"101011111111",
				"101111101111",
				"100110011010",
				"100010001001",
				"110011001110",
				"110111101111",
				"101111101111",
				"100111001110",
				"100010111101",
				"100011001101",
				"101011101111",
				"100111011101",
				"101111101111",
				"110011101111",
				"101010101100",
				"100110101100",
				"100111011111",
				"100011011110",
				"101011011111",
				"101111011111",
				"101111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100011111111",
				"100111111111",
				"100111101110",
				"100111011110",
				"101011101110",
				"101111011110",
				"011110011010",
				"100010101011",
				"100111011110",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011011110",
				"101011101111",
				"101011011111",
				"100011001101",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"101011101111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101011011111",
				"100110111101",
				"011110101100",
				"010110011010",
				"010010011010",
				"011010101011",
				"100111001101",
				"101111101111",
				"110011101111",
				"110011011110",
				"101111011110",
				"100010101011",
				"100010111100",
				"100010111100",
				"100011001101",
				"100011001110",
				"011111001110",
				"011111011110",
				"011111011111",
				"011011011111",
				"011011011111",
				"011011011111",
				"011011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111011110",
				"011011001101",
				"011111001101",
				"011111001100",
				"011110111011",
				"100010111011",
				"100010111011",
				"100010101011",
				"011010001001",
				"011110101011",
				"011110111100",
				"100010111101",
				"100011001110",
				"011111001110",
				"011111001101",
				"011111001110",
				"100011011110",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011111001100",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110111011",
				"010110111100",
				"010110111100",
				"010110111100",
				"010111001100",
				"010111001100",
				"011011001100",
				"011011001100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110101011",
				"011010101011",
				"010110101010",
				"010010011001",
				"001110001000",
				"010010011001",
				"011010011010",
				"100010101011",
				"100010011011",
				"011110001010",
				"011010001001",
				"010110001001",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110101001",
				"010110101001",
				"010110011001",
				"010110101001",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010001001",
				"011010001001",
				"011001111000",
				"010101111000",
				"010101111000",
				"010110001001",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010010101010",
				"010010011010",
				"010010011001",
				"010010011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010110001001",
				"010110011001",
				"010010001000",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011001",
				"011010001001",
				"011010011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"001101111000",
				"001101100111",
				"001101110111",
				"010010001000",
				"010110001001",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001000",
				"010010001000",
				"010001111000",
				"010110001001",
				"011010011010",
				"010110011001",
				"010010001001",
				"010001111000",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010110",
				"011001100110",
				"011001100110",
				"011001110111",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111100",
				"110011001100",
				"110010111100",
				"110011001100",
				"110010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011110",
				"110011011110",
				"110011011101",
				"110011011110",
				"110011011110",
				"101111011101",
				"101111011101",
				"101111011110",
				"101111011101",
				"101111011101",
				"101111011101",
				"110011011110",
				"110011011110",
				"101111001101",
				"101111001101",
				"101111011101",
				"101011001101",
				"101111011110",
				"101011001101",
				"101010111100",
				"100110101011",
				"101111001101",
				"110011011110",
				"101111011110",
				"101111011110",
				"101111001101",
				"100110111100",
				"101111001110",
				"110011011111",
				"101111001110",
				"101111001101",
				"101111011101",
				"101111011101",
				"110011101110",
				"110011011101",
				"100010001000",
				"011110001001",
				"101111011101",
				"101011101110",
				"101011111111",
				"100011101111",
				"101011111111",
				"101111101111",
				"100110011010",
				"011101111000",
				"101010101100",
				"101111001110",
				"100111001101",
				"100010111100",
				"100011001101",
				"101111101111",
				"101011101111",
				"100111011110",
				"110011111111",
				"110011101111",
				"100110101011",
				"100110101100",
				"100111011111",
				"100011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011111111",
				"100111101111",
				"101011111111",
				"100111101110",
				"101111101111",
				"101111011110",
				"110011011110",
				"100010011010",
				"100010011011",
				"100111011110",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100111011111",
				"100111011110",
				"101111101111",
				"101011011110",
				"100111001101",
				"110011101111",
				"101111011111",
				"101111011111",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"100111001110",
				"100010111100",
				"100010101100",
				"011110011011",
				"011010011011",
				"011110111100",
				"011111001101",
				"100011001101",
				"100111011110",
				"100111011110",
				"100111011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"100111001101",
				"011110101011",
				"011010111100",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011110111100",
				"011110101010",
				"100010101011",
				"100110111011",
				"100010101010",
				"011110011010",
				"011110101011",
				"011110111100",
				"011110111101",
				"011111001110",
				"011011001110",
				"011011001110",
				"011111011110",
				"011011001101",
				"011010111101",
				"011010111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011111001100",
				"011010111011",
				"010110111011",
				"011010111100",
				"011011001100",
				"011111001101",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"011010101011",
				"010110001001",
				"010001111000",
				"001110001000",
				"010010001001",
				"010010011001",
				"011010111011",
				"011110111011",
				"100010111100",
				"100010111100",
				"100110111101",
				"100010111100",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010101010",
				"011010101010",
				"011010011001",
				"011010001001",
				"011010011010",
				"011110011010",
				"011110001001",
				"010101111000",
				"010101111001",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010010101010",
				"010110101010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010010001000",
				"010010001001",
				"010110011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"011010011001",
				"011010011010",
				"011110011010",
				"010110001001",
				"010101111001",
				"010001111000",
				"010001111000",
				"001101111000",
				"001101111000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"000100010001",
				"000100100010",
				"001000100011",
				"001100110011",
				"001101000100",
				"010001000100",
				"010001010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001110111",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011110",
				"110011011101",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001101",
				"110011011101",
				"110011011110",
				"101111011101",
				"101111001101",
				"101011001101",
				"101111011101",
				"101111011101",
				"101111001101",
				"101010111100",
				"101010111100",
				"101011001101",
				"101111011101",
				"110011011110",
				"101111011110",
				"101011001101",
				"100110111100",
				"101111011110",
				"110011011111",
				"101111001101",
				"101011001101",
				"101111011101",
				"101111011101",
				"110011011110",
				"101111001101",
				"011101111000",
				"100110101011",
				"101111011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"110011111111",
				"101010111100",
				"100001111000",
				"100110001010",
				"100010011011",
				"100010111100",
				"100111001110",
				"100111011111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101111111111",
				"110011111111",
				"100010011011",
				"100010101100",
				"100111011111",
				"100011101111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110111101111",
				"110011101111",
				"100110011011",
				"100010001001",
				"101010111101",
				"100111011110",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100111101110",
				"101011101111",
				"101011011111",
				"011110011011",
				"100010011010",
				"101010111101",
				"100110011011",
				"100010011011",
				"011110001010",
				"011110011010",
				"011110011011",
				"011110011011",
				"011110011011",
				"011110101100",
				"100010111101",
				"100010111101",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101110",
				"100111101110",
				"101011101111",
				"101011101111",
				"011110111101",
				"011110111100",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011101111",
				"011111011110",
				"011111011110",
				"100011101111",
				"100011101111",
				"100011101110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011011001101",
				"011111001101",
				"100011001100",
				"100010111011",
				"101010111100",
				"101010111100",
				"100110101011",
				"100010011010",
				"100010011011",
				"100010111101",
				"011111001101",
				"011111011110",
				"011011001110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011110101011",
				"100010111101",
				"011110101011",
				"100111001110",
				"100111001110",
				"100110111101",
				"100111001101",
				"100010111100",
				"100010111100",
				"011010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011110101011",
				"011110111100",
				"100011001100",
				"011111001100",
				"011010111011",
				"010110101010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101001",
				"010110101010",
				"010110101010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011010",
				"010110011001",
				"010110001001",
				"011010001001",
				"011110011010",
				"011010001001",
				"010101101000",
				"010101111000",
				"011010001001",
				"011010011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010010101010",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110011001",
				"010010001000",
				"010110001001",
				"010110001001",
				"001101100111",
				"001101100111",
				"010101111000",
				"010110001001",
				"010001111000",
				"010101111001",
				"010001111001",
				"010110001001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110001001",
				"010001111000",
				"010001111000",
				"010110001000",
				"010110001001",
				"010001111000",
				"001101111000",
				"010110011001",
				"011010101010",
				"010110011010",
				"011010101010",
				"010110011001",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"000100010001",
				"000100010010",
				"001100110011",
				"001100110100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101011",
				"101110101011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"110011001100",
				"110011001100",
				"101110111100",
				"101110111011",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111011101",
				"101111001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101010111101",
				"101011001101",
				"101111001101",
				"101111011110",
				"101111011101",
				"101011001100",
				"100110111100",
				"101111001101",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"100010001001",
				"100110101011",
				"101111011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101111111111",
				"101010111011",
				"011001100111",
				"100010001001",
				"100110101100",
				"100111001110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"101011101111",
				"110011111111",
				"100110111100",
				"100010101100",
				"100111011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101111101111",
				"110011101111",
				"101111001101",
				"100010001010",
				"011101111001",
				"101010011011",
				"101111001110",
				"100111011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101110",
				"101111101111",
				"100110111100",
				"011110001010",
				"100110011011",
				"100110001010",
				"100010001010",
				"100010011011",
				"100010101011",
				"100010111100",
				"100010111101",
				"100010111101",
				"100111001110",
				"100111001110",
				"100111011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"011111011110",
				"011111011110",
				"011111101110",
				"011111101111",
				"100011101111",
				"100011011111",
				"101011101111",
				"101011101111",
				"100011001110",
				"011110111101",
				"011110111101",
				"100011001110",
				"011111001110",
				"011111011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111101110",
				"100011101111",
				"011111101110",
				"011111011110",
				"011111001110",
				"100011011110",
				"100111011110",
				"100111001101",
				"101011001101",
				"101010111100",
				"100110011010",
				"100010001001",
				"100010011010",
				"100010011011",
				"100010111100",
				"011110111101",
				"011111011110",
				"011011011110",
				"011011101111",
				"011011011111",
				"011011011110",
				"011111011110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011110111100",
				"100010111100",
				"011110101011",
				"100010011011",
				"100110111100",
				"100110111101",
				"100110111101",
				"100010101100",
				"011110011010",
				"011110011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"010110101011",
				"011010111100",
				"011111001100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"011010011001",
				"011010011010",
				"011010001010",
				"011010001001",
				"010101111000",
				"011010001001",
				"010110001001",
				"010110011010",
				"011010101010",
				"011010101011",
				"010110101010",
				"010110101010",
				"011010111011",
				"010110101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010110001001",
				"010110001001",
				"010101111000",
				"010101111001",
				"011010001001",
				"010101111001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010101111000",
				"011010011010",
				"011110011010",
				"011110101011",
				"011010011010",
				"010110001001",
				"010010001001",
				"010001111000",
				"001101111000",
				"001101111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100011",
				"001100110011",
				"010001000100",
				"010001010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101100110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"101111001101",
				"101111001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111001101",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"100110101011",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111011101",
				"101111011101",
				"110011011101",
				"110011001101",
				"100110011011",
				"101010111100",
				"101011011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101111101111",
				"101010111100",
				"010101010110",
				"011101111000",
				"100110101100",
				"100111011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100111101110",
				"101111111111",
				"101011001110",
				"100010101011",
				"100111011110",
				"100111011110",
				"100111101110",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101111101111",
				"110011111111",
				"110011111111",
				"101111011110",
				"101011001101",
				"100010011010",
				"011001111000",
				"100010001010",
				"110010111101",
				"101111001110",
				"100111011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"101011101111",
				"101011011110",
				"011110001010",
				"011101111001",
				"100110001010",
				"100110011011",
				"100110101100",
				"100110111101",
				"100111001101",
				"100111001110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011011101111",
				"011011101111",
				"011111101111",
				"011111101111",
				"100011011111",
				"100111011111",
				"101011111111",
				"101011101111",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011011110",
				"011111011110",
				"011111001110",
				"100011011110",
				"100111011110",
				"100111001101",
				"101011001101",
				"100110101100",
				"011001111000",
				"011001101000",
				"100110011011",
				"100110101100",
				"100010101100",
				"100010101100",
				"011110111101",
				"011111001110",
				"011011001101",
				"011011011110",
				"011011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011111001101",
				"011011001100",
				"011010111011",
				"011010101011",
				"011110101011",
				"011110101011",
				"011110001010",
				"011001111001",
				"011110001010",
				"011110001010",
				"011110001010",
				"011010001010",
				"011110011011",
				"011010011010",
				"011010011011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"010110101011",
				"010010011010",
				"010010011010",
				"010110101011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010011010",
				"010001111000",
				"001101010111",
				"001101010111",
				"010101111000",
				"010101111001",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001001",
				"011010011010",
				"011010001001",
				"010101111001",
				"011010001001",
				"010101111001",
				"011010011010",
				"010110001001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001001",
				"010001111000",
				"010001111000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010001100111",
				"010001100111",
				"010001111000",
				"010110001001",
				"010110001001",
				"001101100111",
				"001101110111",
				"001101111000",
				"001101111000",
				"010010001000",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101100110",
				"011101100110",
				"011101110110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010011000",
				"100010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111010",
				"101010101010",
				"101010111011",
				"101110111011",
				"101010101010",
				"101010111010",
				"101110111011",
				"101110111011",
				"101110101010",
				"101110101010",
				"101110111010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"110010111011",
				"110011001100",
				"110010111100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"101111001100",
				"101111001100",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"101111011101",
				"101111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"100110101011",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111011101",
				"101111001101",
				"101011001100",
				"110011011101",
				"110011011110",
				"100110101100",
				"101010111101",
				"101011011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101111101111",
				"101111001101",
				"010101010110",
				"011101111000",
				"100110111100",
				"100111011110",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101110",
				"101011111111",
				"101111011110",
				"100010101011",
				"101011011110",
				"101111101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011101111",
				"101111111111",
				"110011111111",
				"110011101111",
				"101111101111",
				"100111001101",
				"100111001101",
				"101011011110",
				"101111011110",
				"100110111100",
				"100110101011",
				"101010111100",
				"101011001101",
				"100111011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"011111101110",
				"011111101110",
				"100111101110",
				"101111101111",
				"100110101100",
				"011101111001",
				"100110011011",
				"101010101101",
				"101010111101",
				"100111001110",
				"100111011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011011101111",
				"011111101111",
				"011111011111",
				"100011101111",
				"100011011111",
				"101011101111",
				"101011101111",
				"100111011111",
				"100011011110",
				"011011001101",
				"011111001110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111011110",
				"100011011110",
				"100011011110",
				"100111011111",
				"100111011111",
				"100010111101",
				"100111001110",
				"100010101100",
				"011010001001",
				"010101101000",
				"010101101000",
				"011110001001",
				"100110101100",
				"100110101100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011111001110",
				"011011001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010111100",
				"010110111011",
				"011011001100",
				"011011001100",
				"011010101011",
				"011110111011",
				"100010111100",
				"100010101011",
				"011010001001",
				"010101101000",
				"011010001001",
				"100010101100",
				"011110011011",
				"011110101100",
				"100010111101",
				"011110111101",
				"011110111100",
				"011110111101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011011001100",
				"011010111100",
				"010110101011",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010111011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101011",
				"010110011001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110001001",
				"011010001010",
				"011010011010",
				"010001111000",
				"010110001001",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"011010001001",
				"011010001001",
				"011010001001",
				"010101111001",
				"010001111000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"001101111000",
				"010001111000",
				"010110001000",
				"011010001001",
				"010101111000",
				"001101010110",
				"000100110100",
				"001101010110",
				"010001111000",
				"010001111000",
				"001101111000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001000100010",
				"001000110011",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011011101",
				"110011011101",
				"110011011101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011011101",
				"101111011101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"100110111011",
				"101010111101",
				"101011001101",
				"101111001101",
				"101111011101",
				"101011001100",
				"101010111011",
				"101111001101",
				"110011011110",
				"101010111100",
				"100110111101",
				"101011011111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"110011101111",
				"110011011101",
				"011001100111",
				"011110001001",
				"101011001101",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100111101110",
				"101011111111",
				"110011101111",
				"100010011011",
				"101011001101",
				"110011101111",
				"101111101111",
				"110011101111",
				"110011111111",
				"110011111111",
				"110011111111",
				"101111101111",
				"100111001110",
				"100010111100",
				"100011001101",
				"100111011110",
				"101111111111",
				"110111111111",
				"110011111111",
				"100110111100",
				"100010101011",
				"100111001101",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011111111",
				"100011111111",
				"100011011110",
				"101111101111",
				"101111001110",
				"100010001010",
				"100010011011",
				"101010111101",
				"101011001110",
				"100111001110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011011111",
				"011010111101",
				"100011011110",
				"100011011111",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111011111",
				"100111011111",
				"101011101111",
				"101011011111",
				"100111001110",
				"100010111101",
				"011110101100",
				"011010011011",
				"011010001010",
				"100010101100",
				"101011011110",
				"101011011110",
				"100110111100",
				"011110101011",
				"011110011011",
				"011110111100",
				"011110101100",
				"011110111101",
				"011110111101",
				"100011001110",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001100",
				"010010111011",
				"010111001100",
				"010111001100",
				"010110111011",
				"011010101011",
				"011110111011",
				"100010101011",
				"011110011010",
				"010110001000",
				"011110011010",
				"100010111100",
				"011010011010",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111101",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111011",
				"011110111100",
				"011010101011",
				"010110101010",
				"010110011010",
				"010010001001",
				"001110001000",
				"001110001001",
				"010110011010",
				"011010101011",
				"011110111100",
				"100010111101",
				"100111001101",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010110011001",
				"010110001001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010101111000",
				"011010011010",
				"011110011010",
				"010101111001",
				"010001100111",
				"010110001001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001110111",
				"011010001001",
				"011001111000",
				"010101100111",
				"001000110101",
				"010001100111",
				"010101111000",
				"010110001001",
				"010001111000",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101100101",
				"010101100110",
				"010101100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011010",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101110111100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001101",
				"110011001100",
				"110011001101",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101111011101",
				"101111011101",
				"101011001100",
				"100110111011",
				"101111001101",
				"101111001110",
				"100110111101",
				"100110111101",
				"101011011111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"110011101111",
				"110111011110",
				"011101111000",
				"100010011010",
				"101011001101",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"101011111111",
				"100111011110",
				"100111101110",
				"101011111111",
				"110011111111",
				"011110011010",
				"100010011010",
				"101111001101",
				"101111011110",
				"110011101111",
				"110111111111",
				"101111011111",
				"100111001101",
				"100010111100",
				"100011001101",
				"100011001101",
				"101011101111",
				"101011111111",
				"101011101110",
				"101011101111",
				"110011111111",
				"101111011110",
				"100110111100",
				"100111001101",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"011111101111",
				"100011111111",
				"100011011101",
				"101111101111",
				"110011101111",
				"100110101100",
				"100010011011",
				"100110111101",
				"100111001110",
				"100011011110",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011101111",
				"100011011111",
				"011111011110",
				"100111101111",
				"100111101111",
				"100011001110",
				"100011001101",
				"100111101111",
				"100111101111",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"100111001101",
				"100010111101",
				"011110101011",
				"011010011011",
				"010110001010",
				"011110111100",
				"100011001101",
				"101011011110",
				"101011011111",
				"101011011110",
				"101111111111",
				"101111101111",
				"100011001101",
				"011010111100",
				"011010101100",
				"011010111101",
				"011111001101",
				"100011001110",
				"011110111101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001110",
				"011111001110",
				"100011001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011011001101",
				"010111001100",
				"010110111100",
				"011010111011",
				"010110101010",
				"011010101010",
				"011110101010",
				"011110101010",
				"010110001000",
				"011010011001",
				"011110101011",
				"010110101011",
				"011010101100",
				"010110101100",
				"010110111101",
				"011011001101",
				"011010111101",
				"011110111101",
				"011110111101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010010101010",
				"010110101010",
				"010110111011",
				"011010111011",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010101011",
				"011010011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"001110001001",
				"010010011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011110111100",
				"100010111100",
				"100011001101",
				"011010101011",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010010011010",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010010001000",
				"010110001001",
				"010110001001",
				"010101111000",
				"011110011010",
				"011110011010",
				"010001101000",
				"001101100111",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010011001",
				"010110011001",
				"010110001000",
				"010001111000",
				"010101111000",
				"010101111000",
				"011001111000",
				"010001010110",
				"010101101000",
				"010101111000",
				"010101111000",
				"010001111000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001010101",
				"010101010101",
				"010101010101",
				"010101010110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010101001",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101110101010",
				"101110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"110011001101",
				"110011001101",
				"101111001101",
				"101111001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101011001100",
				"101111001101",
				"101011001101",
				"101010111100",
				"101010111100",
				"101010111100",
				"101111001101",
				"101111011101",
				"100110111011",
				"100110101011",
				"101111001101",
				"101111001101",
				"101010111101",
				"100010111101",
				"100111001110",
				"100111011111",
				"100111011111",
				"101011101111",
				"101111101111",
				"110011101111",
				"110011011110",
				"100010001001",
				"100110101011",
				"101011001101",
				"100111101111",
				"100111111111",
				"100111111111",
				"101011101111",
				"101011111111",
				"100111101110",
				"100111101110",
				"101011101110",
				"110011101111",
				"100010011010",
				"011001111001",
				"100110101011",
				"101010111101",
				"101010111101",
				"100110111101",
				"100010111100",
				"100010111101",
				"100111011110",
				"101011101111",
				"101011111111",
				"100011011110",
				"101011111111",
				"101011101111",
				"101011101111",
				"110011111111",
				"110011101111",
				"101010111100",
				"100111001101",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100111011110",
				"101111101111",
				"110011011111",
				"101010101100",
				"100110011011",
				"100110111101",
				"100111011110",
				"100111011111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"100011101111",
				"011111011110",
				"011111011110",
				"100111101111",
				"101011101111",
				"101011011111",
				"100011001101",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111001110",
				"100010111101",
				"011010101011",
				"010110011010",
				"010110011010",
				"011010011011",
				"011110111101",
				"100011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111101111",
				"011010111100",
				"010110101100",
				"010110101100",
				"011010111101",
				"011111001110",
				"011011001101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011011001101",
				"011010111100",
				"011110111100",
				"011110111011",
				"011110111011",
				"100010111100",
				"100010111011",
				"010110001000",
				"010110011001",
				"011010011010",
				"011010101011",
				"011111001101",
				"010110111100",
				"011010111101",
				"011011001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"011010111011",
				"010110101011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010010011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010101100",
				"011010101011",
				"100011001101",
				"011111001100",
				"011010101011",
				"010010011010",
				"010010011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110101010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110101001",
				"010110101001",
				"010110101001",
				"010110011001",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010001001",
				"011010001001",
				"011001111001",
				"010001101000",
				"010001111000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011010",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010110001000",
				"010110001000",
				"010110001001",
				"010110001001",
				"010110011001",
				"010010011001",
				"010010011001",
				"010010001000",
				"010010001000",
				"010110001000",
				"011010001000",
				"011001111000",
				"100010001001",
				"011001101000",
				"011001111000",
				"010101100111",
				"010101111000",
				"010110001000",
				"010010001001",
				"010010001001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001000",
				"010001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100100001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000110011",
				"001100110100",
				"010001000100",
				"010001010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110011000",
				"101010011000",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101111001100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101111001100",
				"101111001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"110011001100",
				"101111001100",
				"101111001100",
				"110011001101",
				"101111001101",
				"101111001101",
				"101111001100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001101",
				"101111001101",
				"101010111100",
				"101111001101",
				"101111001101",
				"101011001100",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001100",
				"100010101010",
				"100010101010",
				"101111001101",
				"101111001101",
				"101010111101",
				"100010101100",
				"100111001101",
				"100111011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"101010111100",
				"100010001001",
				"101010111100",
				"101011011111",
				"101011111111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"100111011101",
				"101111101111",
				"101010111101",
				"100010001010",
				"100110011011",
				"100010011011",
				"100110111101",
				"100111001110",
				"101011011110",
				"100111011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"101011101110",
				"110011111111",
				"110011101111",
				"101011001101",
				"100110111100",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011111111",
				"100111101110",
				"101111101111",
				"110011011111",
				"101110111101",
				"100110101100",
				"100110101100",
				"100111001101",
				"100111011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011011110",
				"100011001110",
				"101011101111",
				"101011011110",
				"011110101011",
				"100110111101",
				"101011001110",
				"101011001110",
				"100110111101",
				"100010111100",
				"011110101011",
				"011010011010",
				"010110011010",
				"010010011010",
				"010010011010",
				"011010101100",
				"011111001101",
				"100011001110",
				"100011011110",
				"100011011110",
				"011111011101",
				"011111101111",
				"011111011110",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111101111",
				"011111001110",
				"011010111101",
				"010110111100",
				"011011001101",
				"011010111100",
				"011011001101",
				"011111011101",
				"011011011101",
				"011011011110",
				"011011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011110111100",
				"011110101011",
				"100111001100",
				"100110111100",
				"011110011001",
				"010110001000",
				"011010001001",
				"010110011010",
				"011010101011",
				"011111001101",
				"011010111101",
				"011011001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"011110101011",
				"100010101100",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010111100",
				"011110111100",
				"011010111100",
				"010110111011",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010101011",
				"011010111011",
				"011110111100",
				"011110111100",
				"011010101011",
				"010010001001",
				"010010011001",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101010",
				"010010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010001101000",
				"010001100111",
				"010101111000",
				"010001111000",
				"010110001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010010001000",
				"010010001000",
				"010110001000",
				"010010001000",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"001101110111",
				"010001111000",
				"010110001000",
				"011001111000",
				"011001111000",
				"100010011010",
				"011001111000",
				"010101100111",
				"010001100111",
				"010101111000",
				"010001111000",
				"010001111000",
				"010010001001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000010010",
				"001000100011",
				"001100110011",
				"010001000100",
				"010001000101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"110010111100",
				"101110111100",
				"101110111100",
				"101110111100",
				"101111001100",
				"101111001101",
				"101111001101",
				"101111001100",
				"101110111100",
				"101110111100",
				"101111001101",
				"110011001101",
				"101111001100",
				"101010111100",
				"101111001101",
				"101111001101",
				"101111001100",
				"101010111100",
				"101010111100",
				"101011001100",
				"101011001100",
				"100010101010",
				"100010101010",
				"100110111100",
				"101011001101",
				"101011001110",
				"100010101100",
				"100110111101",
				"101011001110",
				"101011011110",
				"101111101111",
				"101111011110",
				"110111101111",
				"101010111100",
				"100010001010",
				"101011001101",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011101110",
				"110011101111",
				"101111001101",
				"011001101000",
				"100110011011",
				"100110111101",
				"101011001110",
				"101011011111",
				"101011011111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101111101111",
				"110011101111",
				"101011001110",
				"100110111100",
				"100011011110",
				"100011011110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"101011111111",
				"101011011111",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101011011110",
				"101010111100",
				"100110011010",
				"100001111000",
				"100110011010",
				"100010111100",
				"100011011110",
				"100011101111",
				"100011011111",
				"100111011111",
				"100011011111",
				"100011101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011011111",
				"011111011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100111011110",
				"101011011111",
				"011110001010",
				"011001111000",
				"011110011010",
				"011001111001",
				"011001111001",
				"011101111001",
				"100010001011",
				"011110001011",
				"011010101011",
				"011010111101",
				"011011011110",
				"011011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100111101111",
				"100011101111",
				"011011001101",
				"010110111011",
				"011011001100",
				"011111011101",
				"011011001101",
				"011011011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011101",
				"011011011101",
				"011011011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"100110111101",
				"100010101011",
				"010101111000",
				"001101000110",
				"010101111000",
				"100010101100",
				"011110011011",
				"100010111100",
				"011010101100",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101010",
				"011110101011",
				"011010011001",
				"011001111001",
				"010101111000",
				"010101111001",
				"011110011010",
				"010110001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111100",
				"011010111100",
				"010110111100",
				"011010111011",
				"010110101011",
				"011010101011",
				"011110111011",
				"011110101011",
				"011010101011",
				"010010011010",
				"010010001001",
				"011010101011",
				"011010101011",
				"011010101010",
				"010110011010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110111010",
				"010110101010",
				"011010101010",
				"011010101010",
				"011010101010",
				"010110101010",
				"010110011010",
				"010110101010",
				"011010101011",
				"011110101011",
				"011010011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"011010001001",
				"011010001001",
				"011010001001",
				"001101100111",
				"010001111000",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"011010011010",
				"010110001010",
				"010110001001",
				"010110001001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010010011001",
				"010110001001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001000",
				"010101111000",
				"011110011001",
				"011110001001",
				"010101100111",
				"010001010110",
				"010101100111",
				"010101111000",
				"010101111000",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"000100010010",
				"001000100011",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111011",
				"101110111100",
				"101111001100",
				"110011001100",
				"101110111100",
				"101110111100",
				"101010111100",
				"101111001100",
				"110011001101",
				"101111001100",
				"101010111100",
				"101010111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101010111100",
				"101011001100",
				"101011001100",
				"100010101011",
				"100010101011",
				"100110111100",
				"101011001101",
				"101111001110",
				"100110111100",
				"100110111100",
				"101011001101",
				"101111011110",
				"101111011110",
				"101111011110",
				"110011101111",
				"101110111101",
				"100010011011",
				"101011001110",
				"100111011111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011101110",
				"101011011101",
				"101111101111",
				"101111011110",
				"011101111001",
				"100010001011",
				"101011001110",
				"101011011111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101111101111",
				"110011101111",
				"101111011110",
				"100111001101",
				"100011011101",
				"100011011110",
				"100111011111",
				"101011101111",
				"101011111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"100110111101",
				"100110101100",
				"011101111000",
				"011001000110",
				"100001100111",
				"101010111100",
				"100011001100",
				"100011011110",
				"100011101111",
				"100011011111",
				"100111011111",
				"100111011111",
				"100011101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011111",
				"101011101111",
				"100110111100",
				"011101111000",
				"011001111000",
				"011110001001",
				"100010001011",
				"100110011011",
				"100110011100",
				"100110111101",
				"100011001110",
				"011111011110",
				"011011101111",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011101111",
				"011111011110",
				"011111001101",
				"011111001100",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011011110",
				"011111011110",
				"011111011110",
				"100011101111",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011110",
				"011111011101",
				"011011001101",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001100",
				"100011011101",
				"100111011101",
				"100111001101",
				"011110101011",
				"010101111001",
				"010001010111",
				"001101000110",
				"001000110101",
				"011001111001",
				"100010101011",
				"011110011010",
				"100010111101",
				"011010101100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101010",
				"011010101010",
				"011010011010",
				"100010101011",
				"011010001001",
				"010101100111",
				"010101111000",
				"011110011011",
				"011010011010",
				"011010101011",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111011",
				"010110101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101010",
				"011010101010",
				"010110101011",
				"010110111010",
				"011010101010",
				"011010101010",
				"010110101001",
				"010110101010",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"011010011010",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010011010",
				"010001111000",
				"001101101000",
				"010010001001",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010010011001",
				"010010011001",
				"001110011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110001001",
				"011010011001",
				"010101111000",
				"001101010110",
				"001001000101",
				"001101010110",
				"010101110111",
				"010101111000",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000011",
				"010001000100",
				"010101010101",
				"010101100101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111010",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101111001100",
				"101110111100",
				"101010111100",
				"101110111100",
				"101111001100",
				"101111001100",
				"101110111100",
				"101010111100",
				"101010111100",
				"101111001101",
				"101111001100",
				"101010111100",
				"101010111100",
				"101011001100",
				"100110111011",
				"100010101011",
				"100110111100",
				"101011001101",
				"101011001110",
				"100110111101",
				"100110111100",
				"101011001101",
				"101111011110",
				"101011001101",
				"101011011110",
				"101111011110",
				"101111001110",
				"100110101100",
				"100111001110",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011101111",
				"101111111111",
				"101011101110",
				"101111101110",
				"101011011101",
				"101111101110",
				"101111011110",
				"011101111001",
				"011101111010",
				"101011001110",
				"101011011111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"110011101111",
				"101111101111",
				"101011001110",
				"101011011110",
				"100111011110",
				"101011011110",
				"101011011111",
				"101011101111",
				"100111101111",
				"100111111111",
				"101011111111",
				"101011101111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111111111",
				"101011101111",
				"100011001101",
				"011110101100",
				"101011011110",
				"110011011111",
				"101110111100",
				"100010001001",
				"100101111001",
				"101110111100",
				"100011001100",
				"011111011101",
				"100011011111",
				"100011101111",
				"100111101111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100111011110",
				"101111011110",
				"100010011010",
				"011001111000",
				"100010011010",
				"101010101100",
				"101010101101",
				"100110111101",
				"100111001110",
				"100011011111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100111011111",
				"100011011110",
				"011110111100",
				"011110111100",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111011101",
				"100011011101",
				"100011011101",
				"011111001101",
				"100011001101",
				"100011011101",
				"100111011110",
				"011111001101",
				"011010111100",
				"010110011010",
				"011010011010",
				"011110101011",
				"100010101011",
				"011110011011",
				"011010001010",
				"010101111001",
				"100010101100",
				"011110101011",
				"011110111100",
				"011010101011",
				"011010111101",
				"011011001101",
				"010110111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010011010",
				"011110011010",
				"011110011010",
				"011001111001",
				"011001111000",
				"011110011010",
				"011010001001",
				"011010011010",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"011010101011",
				"011010101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110101010",
				"011010111011",
				"011010101010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101011",
				"011010101010",
				"010110011001",
				"010010001000",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101011",
				"011110101011",
				"011010101011",
				"010110011010",
				"010010011001",
				"001110001001",
				"010010001001",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"001110011001",
				"010010011001",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010010001001",
				"010110011001",
				"011010011010",
				"011010011010",
				"010101111000",
				"001101100110",
				"001101010110",
				"010001100111",
				"010001100111",
				"010001110111",
				"010110001000",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100001",
				"001000100010",
				"001100110011",
				"010001000011",
				"010001010100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101110111010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101110111100",
				"101110111100",
				"101110111100",
				"101010111011",
				"101110111100",
				"101111001100",
				"101111001100",
				"101010111011",
				"101010111100",
				"101111001100",
				"101111001100",
				"101010111100",
				"101010111100",
				"101011001100",
				"100110111100",
				"100110101011",
				"100110101011",
				"100110111100",
				"101011001101",
				"101011001101",
				"100110111100",
				"101111001101",
				"101111011110",
				"101011001101",
				"101011011110",
				"101011011110",
				"110011011111",
				"100110111100",
				"100111001101",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111111111",
				"101111101111",
				"101111101110",
				"101011011110",
				"101111101110",
				"110011101111",
				"100010001010",
				"100010001010",
				"101011001110",
				"101011011111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111111111",
				"100111111111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101011001110",
				"101111101111",
				"101111101111",
				"101111011111",
				"101011011110",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011101111",
				"101111101111",
				"110011111111",
				"101011101111",
				"100011001101",
				"011010101011",
				"011110111100",
				"101011011110",
				"101011011111",
				"110011101111",
				"111011111111",
				"110111101111",
				"100110011010",
				"101010101011",
				"100111001101",
				"100011001101",
				"011111011110",
				"100011101111",
				"100111101111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100011101110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011001101",
				"101011011110",
				"101010111100",
				"011110001010",
				"100110011011",
				"100110111101",
				"100111001101",
				"100111001110",
				"100011001110",
				"100011011110",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111101111",
				"011111101111",
				"100011011111",
				"100011011110",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011110",
				"100011011111",
				"100111011111",
				"100011011110",
				"011110111101",
				"011110111101",
				"100011001110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"011110111100",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"011110111100",
				"100011001101",
				"100111001110",
				"101011001110",
				"101011001110",
				"100010101100",
				"011110101011",
				"010110001010",
				"011010111100",
				"011110111101",
				"011010111100",
				"010110111100",
				"011011001101",
				"011010111101",
				"011011001100",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101010",
				"011010011010",
				"011010001001",
				"100010101011",
				"011110001010",
				"011001111000",
				"011010001010",
				"011110011010",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110011001",
				"010110001001",
				"011010011010",
				"011110101011",
				"011010101010",
				"011010101010",
				"011110111011",
				"011110111011",
				"011110111011",
				"011010101010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110011010",
				"010110101010",
				"011010101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"011010111011",
				"011010111011",
				"010010011010",
				"001110001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010101010",
				"010010101010",
				"010010101010",
				"010010011001",
				"010110011001",
				"010110011001",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110011001",
				"011010011010",
				"010110001001",
				"011010001001",
				"011010001001",
				"011010011001",
				"011010001001",
				"010001111000",
				"010001100111",
				"010001111000",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101110111010",
				"101110111010",
				"101010111011",
				"101010111011",
				"101110111011",
				"101110111011",
				"101110111011",
				"101010101011",
				"101010111011",
				"101110111100",
				"101111001100",
				"101010111011",
				"101010111011",
				"101010111100",
				"101111001100",
				"101010111100",
				"101010111100",
				"101010111100",
				"101010111100",
				"100110101011",
				"100110101011",
				"100110111100",
				"100111001101",
				"101011001101",
				"101010111100",
				"101111001101",
				"110011001110",
				"101011001101",
				"100111011110",
				"100111011110",
				"110011101111",
				"100110111101",
				"100011001101",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101110",
				"101111101111",
				"101111011110",
				"110011101111",
				"110111111111",
				"100110011011",
				"100110011011",
				"101011001110",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111111111",
				"100111111111",
				"101011111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011011110",
				"100110101011",
				"101111001101",
				"110011011111",
				"110011011111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101011101111",
				"101111101111",
				"101011011111",
				"100011001101",
				"011010101011",
				"011010111100",
				"100011011110",
				"100111101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011111111",
				"110111111111",
				"101010111100",
				"101010101011",
				"100110111100",
				"100111001110",
				"011111001110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011111111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"100011101110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011101",
				"101011001101",
				"100010011011",
				"100110101100",
				"100110111100",
				"100111001110",
				"100011011110",
				"011111011110",
				"100011101111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011011110",
				"100111011110",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011001101",
				"011010101011",
				"011010011011",
				"011010011011",
				"011010101011",
				"010110101100",
				"011011001101",
				"100011011110",
				"100011011110",
				"011111001101",
				"011110111100",
				"100010111101",
				"100111001101",
				"101011101111",
				"100011001101",
				"010110011010",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110101011",
				"011110101010",
				"100010101100",
				"100110111100",
				"011010001001",
				"010101111000",
				"011010001010",
				"100010101011",
				"011110111100",
				"011010101011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"011010101010",
				"011110101011",
				"100010101011",
				"100010101011",
				"100010101011",
				"100010111011",
				"100010111011",
				"011010101010",
				"010110001001",
				"010001111000",
				"010001111000",
				"010010001001",
				"010110011001",
				"010110011010",
				"010110101011",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010010101010",
				"010110101010",
				"010110101010",
				"010010011001",
				"010010001001",
				"010110001001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010010101010",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010010001001",
				"010010001001",
				"010110011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110010",
				"001100110011",
				"010001000011",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010101010",
				"101010111011",
				"101110111100",
				"101010111100",
				"101010111011",
				"101010111011",
				"101010111100",
				"101010111100",
				"100110111100",
				"101010111100",
				"101110111100",
				"101010101100",
				"100110101011",
				"100110111100",
				"100111001100",
				"101011011101",
				"101010111101",
				"101010111101",
				"101111001101",
				"101011001101",
				"100111011101",
				"100111101110",
				"101111101111",
				"100111001101",
				"100010111100",
				"100111011110",
				"101011011111",
				"101011101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"100110011010",
				"100110101100",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"100111101111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"011001111000",
				"100110011010",
				"101110111101",
				"101111001110",
				"101111001110",
				"101011011111",
				"100111011111",
				"100011001110",
				"011110111100",
				"011110111100",
				"011110111101",
				"011111001101",
				"100011011110",
				"100111101111",
				"100111101111",
				"100111011111",
				"101011101111",
				"101111101111",
				"101011101110",
				"110011101111",
				"110111101111",
				"101111001101",
				"100010011011",
				"100111001101",
				"100011001110",
				"100011011111",
				"011111101111",
				"100011101111",
				"011111101111",
				"100011111111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"101011101110",
				"101011001101",
				"100010011011",
				"100110101100",
				"100010111101",
				"100011011110",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"100111011110",
				"100011001110",
				"011110111100",
				"100111001110",
				"101011001110",
				"101011011110",
				"100111001110",
				"100111001110",
				"100111001110",
				"100111011110",
				"100111011110",
				"011110111101",
				"011010101100",
				"010110011011",
				"010110011010",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"100111011111",
				"100011011110",
				"011010101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001101",
				"011111001100",
				"011010111100",
				"011010111011",
				"011010111100",
				"011110111100",
				"100010111100",
				"100010111100",
				"100010101011",
				"011110011010",
				"010101111000",
				"010101111001",
				"011010001010",
				"011110011011",
				"011110101011",
				"011010101011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110111011",
				"010110111011",
				"010110011010",
				"011010101010",
				"011110101010",
				"010110001001",
				"010001100111",
				"011010001000",
				"011110011010",
				"011010011001",
				"011010011001",
				"010110001001",
				"010110001001",
				"011010101010",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110011010",
				"010010011010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110011010",
				"010010011001",
				"010110011010",
				"011010101010",
				"011010101010",
				"011010101010",
				"011010101011",
				"011010011010",
				"010110011001",
				"010010001001",
				"010010011001",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010011001",
				"101010101001",
				"101010101010",
				"101010101001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101010101011",
				"101010111011",
				"101011001100",
				"100110111011",
				"101010111011",
				"101110111100",
				"101110101100",
				"101010101011",
				"100110111100",
				"100111001100",
				"100111001101",
				"101010111100",
				"100110011011",
				"101110101100",
				"101111001110",
				"100011011101",
				"100011011110",
				"101011101111",
				"101011001110",
				"100010111101",
				"100111001110",
				"101011011110",
				"101011011111",
				"101011011111",
				"101111011111",
				"110011101111",
				"110011101111",
				"110111111111",
				"110011101111",
				"110111101111",
				"110011011110",
				"011110001001",
				"100110101100",
				"101111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101111101111",
				"100010001010",
				"100110011010",
				"101010011011",
				"100110101011",
				"100010101100",
				"011110101100",
				"011110101100",
				"011010101100",
				"100011001101",
				"100011001110",
				"100111011111",
				"100111111111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111011110",
				"101011101111",
				"100111101110",
				"101111101111",
				"110111111111",
				"110011011111",
				"100110011011",
				"100110111101",
				"100011001110",
				"100011011111",
				"011111011111",
				"011111101111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111001101",
				"101011001101",
				"100010011011",
				"100010011011",
				"100110101100",
				"100011001101",
				"100011011110",
				"011111101111",
				"011111101111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011110",
				"011111001101",
				"100011011110",
				"100011011110",
				"011010101011",
				"011110001010",
				"100010011011",
				"100110101100",
				"100010101100",
				"100010101100",
				"011010011011",
				"010110001010",
				"010001111001",
				"010010001001",
				"010010011010",
				"011010101100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111011110",
				"011010111100",
				"011111001101",
				"100011011110",
				"100011011110",
				"011111001101",
				"010110101011",
				"010110101011",
				"011011001101",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011110111100",
				"011110111011",
				"011110101011",
				"010101111001",
				"010001101000",
				"010001100111",
				"011010001010",
				"011010011010",
				"011110011011",
				"011110111100",
				"011110111100",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"010110101011",
				"010110111011",
				"011010101011",
				"011110111011",
				"100010101011",
				"011010001001",
				"010101100111",
				"011001111000",
				"100010101010",
				"011110101010",
				"100010101011",
				"011110101011",
				"011110101011",
				"011110101011",
				"011010101011",
				"010110011010",
				"010110101011",
				"011010101100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010010011010",
				"010010011010",
				"010110011001",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011010",
				"011010101010",
				"011010011010",
				"010110011010",
				"010110001001",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010011010",
				"011010101011",
				"011110101011",
				"011010011010",
				"011010011010",
				"011010011010",
				"010110001010",
				"010010001001",
				"010010001001",
				"010010011010",
				"010110011010",
				"011010101010",
				"010110011010",
				"011010011010",
				"011010011010",
				"010110011001",
				"010110011010",
				"010110001001",
				"010110001001",
				"010110011010",
				"010110001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010100",
				"010101010101",
				"011001100101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100010001000",
				"100110001000",
				"100110011001",
				"101010101001",
				"101010101001",
				"101010101001",
				"100110011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"100110101010",
				"100110111011",
				"101010111100",
				"100110111011",
				"100110101011",
				"101110101100",
				"101110101100",
				"101010101011",
				"100110101011",
				"100110111100",
				"100111001100",
				"100110101011",
				"100010001010",
				"101010101100",
				"101111001110",
				"100011001101",
				"011111011101",
				"101011101110",
				"101011011110",
				"100110111101",
				"100111001101",
				"100111001110",
				"101111101111",
				"101111011111",
				"101111011110",
				"110011101111",
				"110011101111",
				"110011111111",
				"110011101111",
				"110111101111",
				"101111001101",
				"011001111000",
				"100110111100",
				"101011011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"101011101111",
				"100111101111",
				"101011111111",
				"101111101111",
				"101010111100",
				"101110101011",
				"101010101011",
				"101010101100",
				"101010111101",
				"100111001101",
				"100111011110",
				"100111101111",
				"100111011111",
				"101011101111",
				"100111101111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100011011111",
				"100111011110",
				"100111101111",
				"100111101110",
				"101011111111",
				"110011111111",
				"110011101111",
				"101010111100",
				"100110101100",
				"100111001110",
				"100011011111",
				"011111011110",
				"100011101111",
				"011111101111",
				"100011101111",
				"100011011110",
				"100111101111",
				"100111011110",
				"100111011110",
				"100111011111",
				"100111101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111101111",
				"100111011110",
				"100111011110",
				"101011101111",
				"101011101111",
				"101011011110",
				"101011001101",
				"100010011010",
				"011001111001",
				"100010101100",
				"100010111100",
				"100011001110",
				"100011101111",
				"100011101111",
				"011111101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111011111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011111",
				"011111011111",
				"100011011111",
				"011111011110",
				"100011011111",
				"100011011110",
				"011011001101",
				"100011011110",
				"100011011111",
				"011110101100",
				"010101101000",
				"011001101000",
				"011001101000",
				"010101101000",
				"010101111001",
				"011010001010",
				"011010101011",
				"011010101100",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111011110",
				"100011001110",
				"011010111100",
				"010110011011",
				"010110101011",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011111001100",
				"011010101011",
				"010110011010",
				"010110001001",
				"011010011010",
				"010101111001",
				"010001111000",
				"011010011010",
				"011010011010",
				"011110101011",
				"011110111100",
				"011010101011",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110101010",
				"011010011010",
				"011110101011",
				"100010011010",
				"011110001001",
				"011110001001",
				"100110101011",
				"100010101011",
				"011110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010010101010",
				"010010101010",
				"010010011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010110011001",
				"010110011010",
				"011010101010",
				"011010011010",
				"011010011010",
				"011110101011",
				"011010011010",
				"011110011010",
				"011110011011",
				"011110011011",
				"011110101011",
				"011110101011",
				"011010011010",
				"010110001001",
				"010001111001",
				"010001111001",
				"010010001001",
				"010110011010",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110001001",
				"010110011001",
				"010110011010",
				"010010001001",
				"010010001001",
				"010110011001",
				"011010011010",
				"011010001010",
				"010110001001",
				"010001111001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110010",
				"001100110011",
				"010001000100",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"101010011001",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110101010",
				"101010101010",
				"101010111011",
				"100110101010",
				"101010111011",
				"101010111011",
				"101010111011",
				"101110101011",
				"101110101011",
				"101110101011",
				"100110101011",
				"100110111100",
				"100111001100",
				"101010101100",
				"100010001001",
				"101010011011",
				"101010111101",
				"100111011110",
				"011111011101",
				"100111101110",
				"101111101111",
				"101011001101",
				"100110111101",
				"101011011110",
				"101011011111",
				"101011001110",
				"110011011111",
				"110011101111",
				"110011111111",
				"101111101111",
				"101011011110",
				"110111101111",
				"110111011111",
				"100010011010",
				"101011001101",
				"101011011110",
				"100111011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111001101",
				"100010001001",
				"100110001010",
				"101010101100",
				"100110111101",
				"101011011110",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011101110",
				"100111101111",
				"101011111111",
				"101011101111",
				"110011101111",
				"110011001110",
				"100110101100",
				"100111001110",
				"100011011110",
				"011111011110",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111011110",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011101111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111101111",
				"101011101111",
				"100111011110",
				"100111001110",
				"100010111100",
				"011010001010",
				"010101101000",
				"010101010111",
				"100010001010",
				"100110111101",
				"011110111100",
				"100111101111",
				"100011101111",
				"011111011110",
				"100011101111",
				"100011101111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"011111011111",
				"011111101111",
				"100011101111",
				"011111101111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"100111011110",
				"100010001010",
				"011001010111",
				"011001101000",
				"100010011011",
				"011110011011",
				"100010111101",
				"011110111101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011011011110",
				"011011001110",
				"011011001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001110",
				"011111001110",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"100011011110",
				"011110111100",
				"010110011010",
				"011010111100",
				"011111001101",
				"011010111100",
				"011111001101",
				"011111001101",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011001101",
				"011111001100",
				"010110101011",
				"010010001001",
				"010010001001",
				"011010101011",
				"100011001101",
				"100111001101",
				"100111001101",
				"100010111100",
				"010110001010",
				"010110001001",
				"011010101011",
				"011110111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110111100",
				"010110111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"010110111011",
				"010110101011",
				"011010111011",
				"010110011010",
				"011010011010",
				"100010101011",
				"100110011010",
				"100010001001",
				"100010001001",
				"100110101011",
				"011010101010",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011110011010",
				"010101111001",
				"010101111001",
				"010101111001",
				"011010001010",
				"010101111000",
				"010101111001",
				"010110001001",
				"010110011010",
				"011010011010",
				"011010011011",
				"011010101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010011001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110011010",
				"010010001001",
				"010010001001",
				"010001111001",
				"010010001001",
				"010010001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010000110011",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011001100110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110101001",
				"100110011001",
				"100110011001",
				"101010101001",
				"101010101001",
				"100110101001",
				"100110101001",
				"101010101010",
				"101010101010",
				"100110101010",
				"100110101010",
				"100110111011",
				"101010101011",
				"101110101011",
				"101110101011",
				"101010101011",
				"101010101011",
				"100110111011",
				"100111001100",
				"101010111100",
				"100110011010",
				"101010011011",
				"101010111100",
				"100111011101",
				"100011011101",
				"100111101110",
				"101111101111",
				"101010111101",
				"101010111101",
				"101011011110",
				"101011011110",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111101111",
				"101011011110",
				"101011011110",
				"110111101111",
				"111011101111",
				"100110101011",
				"100110111100",
				"101011011110",
				"100111011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"110011011101",
				"011101111000",
				"011101111000",
				"101010111100",
				"101111011110",
				"100111011110",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100111101111",
				"100111101111",
				"100011101110",
				"100111111111",
				"100111111111",
				"100111101110",
				"101111101111",
				"110011011111",
				"100110101100",
				"101011001101",
				"100111011110",
				"100011011111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111011110",
				"100010111101",
				"100010111101",
				"100111001110",
				"101011001110",
				"100110101100",
				"100010001010",
				"011001011000",
				"100110001011",
				"100010101100",
				"011110111100",
				"100011011110",
				"011111011110",
				"100111101111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111101111",
				"011111101111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111001101",
				"100111011101",
				"101110111101",
				"011101101000",
				"011001101000",
				"100010011011",
				"100010101100",
				"100010111101",
				"011110111100",
				"100011001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011011001110",
				"011011001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011110111101",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"100011011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"011010111100",
				"010110011010",
				"010010001001",
				"010010011010",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011110111100",
				"100011001101",
				"100111011110",
				"100011001101",
				"011010011010",
				"010110001001",
				"011010011011",
				"011110111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"011010111011",
				"011011001100",
				"011110111100",
				"011010101011",
				"011110011010",
				"100110101011",
				"100010011010",
				"011101111001",
				"011110001001",
				"100010101010",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"011010011010",
				"011110101011",
				"011010011010",
				"010001101000",
				"001101010110",
				"010101111000",
				"011010001001",
				"011010011010",
				"010110001010",
				"011010011010",
				"011010011011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010010011010",
				"010010011010",
				"010110011010",
				"010010011010",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110011010",
				"010110001001",
				"010110001010",
				"010010001001",
				"010110001010",
				"010110011010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010101010100",
				"010101010101",
				"011001100101",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101001",
				"100110011010",
				"100110101010",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010101011",
				"100110111011",
				"100110111100",
				"101010111100",
				"101010101011",
				"100110011010",
				"101010101100",
				"100111001101",
				"100011011101",
				"100111011110",
				"101111101111",
				"101111001101",
				"101010111101",
				"101011001110",
				"101011011110",
				"110011011111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101011011111",
				"110011011111",
				"111011101111",
				"101010111101",
				"100010111100",
				"101011011111",
				"100111011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"110011011110",
				"011101111000",
				"010101100111",
				"100110111100",
				"101111101111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111011111",
				"100111011111",
				"100011011111",
				"100111101111",
				"100111111111",
				"100011101111",
				"100111101110",
				"101111101111",
				"110011011111",
				"101010111101",
				"101011001101",
				"101011011110",
				"101011101111",
				"101011101111",
				"100111011110",
				"101011011111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011011111",
				"100111011110",
				"100011001101",
				"100010111101",
				"100010111101",
				"100111001110",
				"101111011111",
				"110011101111",
				"110011101111",
				"110111011111",
				"101010001011",
				"100001111001",
				"100110111101",
				"011110111100",
				"011111001101",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"011111101111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011111",
				"011111101111",
				"011111011110",
				"011111011110",
				"100011101110",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111001101",
				"100011001101",
				"101111001101",
				"100010011010",
				"011110001010",
				"100010111100",
				"100010111100",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101100",
				"011110111100",
				"100111001110",
				"100011001101",
				"100010111100",
				"100111001101",
				"100011001101",
				"100111001110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011110111100",
				"011010011011",
				"010110011010",
				"010010011010",
				"010010011010",
				"010110101011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111101",
				"100011001101",
				"011110111100",
				"011111001101",
				"100011001101",
				"100011001101",
				"011110111100",
				"010110101011",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"010110111100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"100010101011",
				"100010011010",
				"011110001001",
				"011110001001",
				"100010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010010011001",
				"010010011001",
				"010110011010",
				"010110011010",
				"011110101011",
				"011010001001",
				"001101010111",
				"010101111000",
				"011010001010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010011010",
				"010010011010",
				"010010011001",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001010",
				"010110011010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001000100010",
				"010000110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010001000",
				"100010000111",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110101010",
				"101010101010",
				"101010011010",
				"101010011010",
				"101010101010",
				"100110101010",
				"100110101011",
				"100110111011",
				"101010111011",
				"101110111100",
				"100110011010",
				"100110101011",
				"100111001100",
				"100111011101",
				"100111001101",
				"101011011110",
				"110011001110",
				"101110111101",
				"101111001101",
				"110011101111",
				"110011101111",
				"101111011110",
				"101011011110",
				"100111001110",
				"101011101111",
				"101111101111",
				"101111011111",
				"110111101111",
				"101111011110",
				"100010111100",
				"100111011110",
				"100111011110",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110111101111",
				"100110011010",
				"011001101000",
				"100110101100",
				"101111011111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"101011101111",
				"101111101111",
				"101111001110",
				"101010111101",
				"101010111101",
				"101011011111",
				"101111101111",
				"101111011111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111111111",
				"101111111111",
				"101111101111",
				"101011011111",
				"100111011110",
				"100011001110",
				"011110111101",
				"011110111101",
				"100011001101",
				"100111011110",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110111101111",
				"110011001110",
				"100010001010",
				"100010111100",
				"011110111100",
				"011111001101",
				"100011011111",
				"011111001110",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"011111101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011111",
				"100011101111",
				"100011011110",
				"100011011110",
				"011111011101",
				"011111001101",
				"011111001100",
				"011111001100",
				"100011001100",
				"101011001101",
				"100110101011",
				"100010101011",
				"100010111100",
				"011111001100",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011110111011",
				"011110101011",
				"100010111101",
				"100111001101",
				"100111001101",
				"101011001110",
				"100111001101",
				"100111001101",
				"100011001101",
				"011111001101",
				"011010111100",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010111011",
				"011010111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"011110111100",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011110111100",
				"011110101011",
				"011010001001",
				"010101111000",
				"011001111001",
				"011110011010",
				"011110011010",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"011010111100",
				"011010111100",
				"010110101100",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010011010",
				"010010101010",
				"010110101010",
				"010110011010",
				"011010101010",
				"011110011011",
				"011010001001",
				"011010001001",
				"010110001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010010011001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"010110001001",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010010",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100110",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110001000",
				"100010000111",
				"100010000111",
				"100110011000",
				"100110011000",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010011010",
				"100110101010",
				"101010101010",
				"101010101011",
				"101010101011",
				"101010111100",
				"100110011010",
				"100110101011",
				"100110111100",
				"100111001101",
				"100111001101",
				"101011001101",
				"110011011110",
				"101010111100",
				"101010111100",
				"110111101111",
				"101111011110",
				"101011011110",
				"101011011110",
				"100111001110",
				"101111101111",
				"101111101111",
				"101111011110",
				"110011101111",
				"101111101111",
				"100010111100",
				"100111001110",
				"100111011110",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110111101111",
				"101010101011",
				"011110001001",
				"101010111101",
				"101111011111",
				"100111101111",
				"100111111111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101111011111",
				"100010011011",
				"011110001010",
				"100110101100",
				"101011001110",
				"101111001110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101011011111",
				"100111011110",
				"100011001101",
				"011110111100",
				"011110101100",
				"011110111101",
				"100011001110",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011011111",
				"101011011111",
				"101111011111",
				"110011101111",
				"101010111101",
				"011010011010",
				"011110111100",
				"100111011110",
				"011111001101",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011110",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011011110",
				"100011001101",
				"100011011101",
				"100011001101",
				"100011001101",
				"100111011101",
				"101011011101",
				"101010111101",
				"011110011010",
				"011010001001",
				"011110111011",
				"011111001101",
				"011011001101",
				"011011001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111001110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001101",
				"011110111100",
				"011010011010",
				"010001111000",
				"011010001001",
				"100010101011",
				"100010101011",
				"100010101011",
				"011010001010",
				"010110011010",
				"010110011010",
				"010010011010",
				"010010011010",
				"010010011010",
				"010110101011",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011111001101",
				"011111001101",
				"011011001100",
				"011010111100",
				"011111001101",
				"100011001101",
				"011110111100",
				"010110011010",
				"010110101010",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101011",
				"010110001001",
				"010001101000",
				"010101111000",
				"011010001001",
				"011110011010",
				"011010011010",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010010101010",
				"010110101010",
				"010110101010",
				"010110011001",
				"011110011010",
				"011010001010",
				"010101111001",
				"010001111000",
				"010110011010",
				"010110101010",
				"010110011010",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010010101010",
				"010010101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001001",
				"010010001000",
				"010010001000",
				"010110001001",
				"010110001001",
				"010110001000",
				"010101111000",
				"010101100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000001",
				"000100010001",
				"001000100010",
				"001000100010",
				"001100110011",
				"010001000100",
				"010001000100",
				"010101010101",
				"010101010101",
				"011001100101",
				"011001100110",
				"011101110111",
				"011101110111",
				"011101110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100110001000",
				"100110001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101011",
				"101010101011",
				"100110101010",
				"100110101011",
				"100110111100",
				"101011001101",
				"101011001101",
				"101011001101",
				"110011011110",
				"101010111100",
				"101010101011",
				"110011001101",
				"101011001101",
				"100111011110",
				"100111011111",
				"100111011110",
				"101111011111",
				"101111011111",
				"101011011111",
				"110011101111",
				"110011101111",
				"100010111100",
				"100011001101",
				"100111011110",
				"101011011111",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110011001101",
				"011101111001",
				"011101111001",
				"101111001110",
				"101111011111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101111101111",
				"100110011011",
				"011001101000",
				"011110001010",
				"100010011011",
				"100110011011",
				"100010101100",
				"100010101100",
				"100010101100",
				"011110101100",
				"011110111100",
				"100010111101",
				"100010111101",
				"100011001110",
				"100111011111",
				"100111101111",
				"100111111111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"100010101100",
				"011010011011",
				"100011001101",
				"100011001110",
				"100011101111",
				"011111011111",
				"011111101111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"101011011110",
				"101011011110",
				"100111001101",
				"100111001100",
				"100010101011",
				"011001111000",
				"011001111000",
				"011010001001",
				"011110101011",
				"100011001101",
				"011011001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011011001101",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010011010",
				"001001010110",
				"001101010110",
				"010101111000",
				"011010001001",
				"011110011010",
				"011010001001",
				"011010011010",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011111001100",
				"011010111100",
				"011110111100",
				"011110111100",
				"100010111101",
				"100010111101",
				"011010101011",
				"010110011010",
				"010010001001",
				"010110011010",
				"011110101100",
				"100010101100",
				"011110001010",
				"010101111000",
				"010110001001",
				"011110101011",
				"011010101011",
				"010110101010",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110011010",
				"011010011001",
				"100010011011",
				"011110001010",
				"010101111000",
				"010101111000",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"011010011001",
				"011010001001",
				"011010001000",
				"010101100111",
				"010101100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001000100010",
				"001000100010",
				"001100110011",
				"001100110011",
				"010001000100",
				"010101010101",
				"011001100101",
				"011001100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010001000",
				"100010001000",
				"100010001000",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010001000",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011010",
				"101010101010",
				"101010101011",
				"100110101011",
				"100110101011",
				"100110101011",
				"100110111100",
				"101010111100",
				"101011001101",
				"101011001101",
				"101111001101",
				"101111001101",
				"101010011010",
				"100110001010",
				"100110111100",
				"100111011101",
				"100111011110",
				"100111011111",
				"101111011111",
				"101011001111",
				"101011011111",
				"101111101111",
				"110011101111",
				"101011001101",
				"100010111101",
				"100111011110",
				"101011011111",
				"100111011111",
				"101011011111",
				"101111101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"110111101111",
				"101110111100",
				"011001010111",
				"011101111001",
				"101111001110",
				"101111011111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011111111",
				"100011101111",
				"100111101111",
				"101111101111",
				"101110111110",
				"011101101001",
				"100001111001",
				"100010001010",
				"100010001010",
				"100010011011",
				"100010011100",
				"100010101100",
				"100111001101",
				"100111001110",
				"101011011111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100011101111",
				"011111011110",
				"011111101111",
				"100011101111",
				"100011111111",
				"011111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"101011101111",
				"101011101111",
				"101111011111",
				"011010011011",
				"011110111100",
				"100011011111",
				"011111011110",
				"011111101111",
				"011111101111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100111011111",
				"100011101111",
				"100011101110",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111001110",
				"100111001101",
				"100110111100",
				"100010101011",
				"011110011001",
				"010001010110",
				"001100110101",
				"011001111000",
				"100010011011",
				"100010111100",
				"100011001101",
				"011111001101",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011011001100",
				"011010111100",
				"100011001100",
				"100011001100",
				"011010001001",
				"010001100111",
				"011001111001",
				"011110001010",
				"100010011011",
				"100110111100",
				"100010111100",
				"011110111100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001101",
				"011111001100",
				"010110101011",
				"010110101010",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010111011",
				"011111001100",
				"100011001101",
				"011110111100",
				"011010101011",
				"011010011011",
				"010110011011",
				"010110011010",
				"011110111100",
				"011010101011",
				"011110101011",
				"100110111100",
				"100111001101",
				"100010101100",
				"010110001001",
				"001101111000",
				"010110011010",
				"010110011010",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110101100",
				"011010101011",
				"011010101011",
				"010110101010",
				"011010101011",
				"011010011010",
				"011110011010",
				"100010011010",
				"011101111001",
				"011001111001",
				"010101111001",
				"011010011010",
				"011010101010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011000",
				"010110001000",
				"011110011001",
				"011110011001",
				"011110011001",
				"011001110111",
				"010101100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100010001",
				"001000100010",
				"001100110010",
				"010001000011",
				"010001000100",
				"010101010101",
				"011001010101",
				"011001100110",
				"011101110110",
				"011101110111",
				"011101110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100110001000",
				"100110001000",
				"100110001000",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101011",
				"100110101010",
				"101010101011",
				"100110101010",
				"100110101011",
				"101010111100",
				"101010111101",
				"101011001101",
				"101011001101",
				"110011011110",
				"101010011011",
				"011001100111",
				"100110111100",
				"100111001101",
				"100011011110",
				"100111011111",
				"101111011111",
				"101011001110",
				"101011011111",
				"101011101111",
				"110011101111",
				"101111011111",
				"100010111100",
				"100111011110",
				"101011011111",
				"101011001110",
				"101011011111",
				"101111101111",
				"101011011111",
				"101011011111",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110111101111",
				"110011001110",
				"011001101000",
				"100010001010",
				"110011001111",
				"101011011111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100011111111",
				"100011111111",
				"100111101111",
				"101111101111",
				"110011001110",
				"011101101000",
				"011101101001",
				"011101111001",
				"100010001010",
				"100110101100",
				"101011001110",
				"101011011110",
				"101011101111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100011101111",
				"011111101111",
				"011111101111",
				"011111101111",
				"011111101110",
				"011111101110",
				"100011111111",
				"100011111111",
				"100011101111",
				"100011101110",
				"101011101111",
				"101111101111",
				"100010111101",
				"100010111101",
				"100011001101",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011101111",
				"100011011111",
				"100111011111",
				"100111101111",
				"100111101111",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001110",
				"100111011110",
				"100011001101",
				"100010111100",
				"011110101011",
				"100010111011",
				"100010101011",
				"010101111000",
				"011001100111",
				"011101111001",
				"100010011011",
				"100010111100",
				"100011001110",
				"011011001101",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011011001110",
				"011111011110",
				"011111011110",
				"011011011110",
				"011011011110",
				"011011011110",
				"011111011101",
				"011111011101",
				"011111001101",
				"011111001101",
				"011111011101",
				"011111011110",
				"011111011101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011010111100",
				"011110111011",
				"100111001100",
				"100010101011",
				"010101111000",
				"011010001001",
				"100010011011",
				"011110011011",
				"100010101100",
				"011110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011011001101",
				"011010111100",
				"010110111100",
				"011010111100",
				"011011001100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011111001101",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"100010111100",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010101011",
				"010110011010",
				"010110001001",
				"010110011010",
				"011010101011",
				"011010101100",
				"011010101011",
				"011010101100",
				"011110101011",
				"011110101011",
				"100010111100",
				"100111001101",
				"011110111100",
				"010110011010",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010101011",
				"011010101011",
				"011010101100",
				"011010101100",
				"011110111100",
				"011110111100",
				"011110101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011110101011",
				"010101111000",
				"010001010110",
				"011110001001",
				"011001111001",
				"010101111001",
				"011010011010",
				"011010011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011001",
				"010110011001",
				"010110011000",
				"010110001000",
				"011110011001",
				"011110011001",
				"100010011001",
				"011101110111",
				"011001100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"010001000011",
				"010101010100",
				"010101010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"100110011000",
				"100110011001",
				"101010101010",
				"101010101010",
				"100110011010",
				"101010101011",
				"101010101011",
				"101010101011",
				"101010111100",
				"101111011110",
				"100110111100",
				"101111001101",
				"101111001101",
				"011001111000",
				"011110011010",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101011011111",
				"101111101111",
				"110011101111",
				"100010111101",
				"100111001110",
				"101011011110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111101111",
				"101111011111",
				"101111101111",
				"101111101111",
				"110011111111",
				"101111101111",
				"101011011110",
				"101011001101",
				"101111011110",
				"110111101111",
				"111011111111",
				"011110001010",
				"100001111010",
				"101111001110",
				"101011011110",
				"100111101111",
				"100011101111",
				"100111111111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101011111111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111111111",
				"100111101111",
				"101011011110",
				"110011011111",
				"100010001010",
				"010001000110",
				"011001010111",
				"101010101100",
				"100110101100",
				"100111001110",
				"100011001110",
				"100011011110",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100011101110",
				"101011101111",
				"101111101111",
				"100110111101",
				"100010111101",
				"101111011111",
				"100111011110",
				"100011011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100111011111",
				"100111011111",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011001101",
				"011010111100",
				"011010101011",
				"011010101011",
				"100011001101",
				"101011011110",
				"101011101111",
				"101111011111",
				"100110101100",
				"011101111010",
				"011010001010",
				"011110101100",
				"011110111100",
				"011111001101",
				"100011011111",
				"011011001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111011110",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111011",
				"011110111011",
				"100111001100",
				"011010001001",
				"011001111001",
				"011010001010",
				"011010011011",
				"100011001101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011010111100",
				"010110101011",
				"011010101010",
				"100010111100",
				"100010111100",
				"011110011011",
				"100010111100",
				"011110111100",
				"100011001101",
				"100011001110",
				"100011001101",
				"100011001101",
				"011110111101",
				"011010111100",
				"010110011010",
				"010010011010",
				"010110011010",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010011010",
				"010110001001",
				"010110011010",
				"011010101011",
				"010110011010",
				"010110101010",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011010101011",
				"010110001010",
				"010001100111",
				"001101010111",
				"010101111001",
				"011010001001",
				"010110001001",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101010",
				"011010101010",
				"010110011010",
				"010110011001",
				"010110011001",
				"011010011001",
				"011010011001",
				"011110011001",
				"100110101010",
				"100110011010",
				"011101110111",
				"011001100111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"001000010001",
				"001000100010",
				"001100110010",
				"010001000011",
				"010001000100",
				"010101010100",
				"011001010101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100001110111",
				"100001110111",
				"100001110111",
				"100010000111",
				"100010000111",
				"100010000111",
				"100110001000",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101010",
				"100110011010",
				"101010101011",
				"101010111100",
				"101010111100",
				"101111001101",
				"101010111100",
				"101011001101",
				"101111001101",
				"100010011010",
				"011110011010",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101011011111",
				"101111011111",
				"101111101111",
				"101011011110",
				"100111001101",
				"101111011110",
				"101111011110",
				"101011001101",
				"101111011110",
				"110011101111",
				"110011101111",
				"101111101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"110111111111",
				"101010111101",
				"100010001010",
				"101010111101",
				"100111001110",
				"100111101111",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011111111",
				"101111101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101110",
				"100111011110",
				"110011101111",
				"100110101011",
				"010101000110",
				"010101010111",
				"100110011011",
				"100110111101",
				"101011011111",
				"100111101111",
				"100011011110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011101110",
				"100111101111",
				"101011101111",
				"101011001111",
				"101010111110",
				"101111011111",
				"101011011110",
				"100111011110",
				"100011011110",
				"100011011110",
				"100011011111",
				"100011001111",
				"100011001110",
				"100111011110",
				"100111011110",
				"101011011111",
				"100111011110",
				"100111001110",
				"100111011110",
				"100111011111",
				"100111011110",
				"011110111100",
				"010110011011",
				"010110101011",
				"011010101100",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011111",
				"101011101111",
				"101011001110",
				"011110011011",
				"011010001010",
				"011110101100",
				"011110111101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111011101",
				"011111011101",
				"011111011101",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"100011001100",
				"011110101010",
				"100111001100",
				"011110011010",
				"010101111001",
				"011010001010",
				"011110111101",
				"011110111101",
				"011011001101",
				"011111001110",
				"011111001110",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011110111100",
				"011010111100",
				"011111001100",
				"011010111011",
				"010110001001",
				"011110011010",
				"101011001101",
				"100110111100",
				"100111001101",
				"100010111101",
				"011110111100",
				"011010101011",
				"011010011011",
				"011010011011",
				"010110011011",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"100011001101",
				"011010101011",
				"010110011001",
				"010010011010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110111011",
				"010110111100",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011110101011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010101011",
				"011010011011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010011010",
				"010001101000",
				"010001101000",
				"011010011010",
				"011010011010",
				"010110011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"011010101010",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010011001",
				"011010011001",
				"011110011010",
				"100010101010",
				"100110101010",
				"100010011001",
				"011001110111",
				"011101110111",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"001000010001",
				"001000100010",
				"001100110011",
				"010001000011",
				"010001000100",
				"010101000100",
				"010101010100",
				"010101010101",
				"011001010101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110110",
				"011101110110",
				"011101110110",
				"011101110110",
				"100001110111",
				"100010000111",
				"100010000111",
				"100110011000",
				"100110011000",
				"100110011000",
				"100110011001",
				"101010101010",
				"101010101010",
				"100010001001",
				"100110011001",
				"101010101011",
				"101010111100",
				"101010111100",
				"101111001101",
				"101010111100",
				"101111001101",
				"101010111100",
				"011110001001",
				"101010111100",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011111",
				"101111011111",
				"101111011111",
				"101011001101",
				"110011011111",
				"110011011110",
				"101111001101",
				"110011011111",
				"110011101111",
				"101111101111",
				"101011011110",
				"100111011110",
				"100111011110",
				"101011011111",
				"101011101111",
				"101111101111",
				"101111011111",
				"101111011110",
				"110011111111",
				"110011101111",
				"100010001010",
				"100110101100",
				"100111011110",
				"100011101110",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"101011011111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011011110",
				"110011101111",
				"101110111101",
				"011001010111",
				"011001010111",
				"100010001010",
				"101010111101",
				"100111011110",
				"100011011110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101110",
				"100011101110",
				"100111101111",
				"101011011111",
				"101011001111",
				"101010111110",
				"101010111101",
				"101111011111",
				"101011011110",
				"100011011110",
				"100011001110",
				"100111011111",
				"101011011111",
				"101011011111",
				"101011101111",
				"101011101111",
				"100111011111",
				"100111011111",
				"100111011110",
				"011110111101",
				"011010101011",
				"010110011011",
				"011010101100",
				"011111001101",
				"011111001110",
				"100011011110",
				"100011011111",
				"100111011111",
				"100011011110",
				"100011001110",
				"100011001110",
				"100011001110",
				"101111011111",
				"100111001110",
				"011110011100",
				"011010101011",
				"011110111101",
				"011111001101",
				"011011001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011110111100",
				"100010111100",
				"100110111100",
				"100010101011",
				"011001111000",
				"011001111001",
				"011110011011",
				"100010111101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011111001101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011111001100",
				"011010111100",
				"011010111011",
				"011111001100",
				"011110111011",
				"010001111000",
				"010001100111",
				"011010001001",
				"011110011010",
				"011010011011",
				"011010011011",
				"010110011011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011011",
				"010110101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"100010111100",
				"010110101010",
				"010010011001",
				"010110011010",
				"010110101010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110111011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"011010101011",
				"011110101100",
				"011110111100",
				"100010111100",
				"011110101100",
				"010110001001",
				"001101101000",
				"010110001001",
				"010110001001",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"011010111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101010",
				"010110101010",
				"010110101010",
				"011010101010",
				"011010011001",
				"011110101010",
				"100110111011",
				"100110101011",
				"011001111000",
				"010001010101",
				"011001100110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"000100010001",
				"001000010001",
				"001000100010",
				"001100100010",
				"001100110010",
				"001100110011",
				"010000110011",
				"010001000011",
				"010101010100",
				"010101010101",
				"011001010101",
				"011001100101",
				"011101100110",
				"011101100110",
				"011101110110",
				"011101110110",
				"011101110111",
				"100010000111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101011",
				"100110011001",
				"100110011001",
				"101010101011",
				"101010111100",
				"101010111011",
				"101010111100",
				"101010111011",
				"101110111100",
				"101010111100",
				"100010011010",
				"100010101011",
				"101011001101",
				"101011011101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011111",
				"101111011110",
				"101010111101",
				"101011001101",
				"110011011111",
				"110111101111",
				"110111101111",
				"110011011111",
				"101011011110",
				"100111001101",
				"100111011110",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011011110",
				"101111101111",
				"101111101111",
				"110011101111",
				"110011101111",
				"100110011011",
				"100110011011",
				"101011011110",
				"100011011110",
				"100011101111",
				"100011101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111011111",
				"101011011111",
				"101111101111",
				"101111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101110",
				"110011011110",
				"101110111100",
				"011101100111",
				"011001010111",
				"100010011010",
				"101111001110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011101110",
				"100011101110",
				"100111101111",
				"100111011111",
				"101011011111",
				"100110111101",
				"011110011010",
				"100010101011",
				"101011011110",
				"100111011110",
				"100111001110",
				"101011011111",
				"101011011111",
				"100111001110",
				"100111001110",
				"100111001110",
				"100011001101",
				"011010101100",
				"010110011011",
				"011010101100",
				"011110111101",
				"011111001110",
				"011111001110",
				"011111001110",
				"100111101111",
				"100011011111",
				"100011011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"101011011111",
				"101011011111",
				"100111001110",
				"011010111100",
				"011010111100",
				"011010111101",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011101",
				"011111001101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110101010",
				"011110011010",
				"010101101000",
				"010001010111",
				"011001111010",
				"011110011011",
				"100010111101",
				"011010111101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011010111101",
				"011011001100",
				"011011001100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001100",
				"011111001100",
				"011110101011",
				"001101010110",
				"001001000101",
				"010110001001",
				"010001111001",
				"010110001010",
				"010110011010",
				"011010101011",
				"011110101100",
				"011110101100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010101011",
				"011110111100",
				"011110111100",
				"010110011010",
				"010110011010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101011",
				"011010111011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011110111100",
				"011010101011",
				"011110111100",
				"011010111100",
				"011010101011",
				"010110101011",
				"010010011010",
				"010010011010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011010011010",
				"010010001001",
				"010001111000",
				"010110011010",
				"010110101010",
				"010110101010",
				"010110101010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010011010",
				"011010011010",
				"100010101011",
				"100010111011",
				"100010101010",
				"011010001000",
				"010101100110",
				"010101010110",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000000",
				"000100010000",
				"000100010001",
				"001000100010",
				"001100110010",
				"010000110011",
				"010001000100",
				"010101000100",
				"011001010101",
				"011001100101",
				"011001100101",
				"011001100101",
				"011001100110",
				"011101100110",
				"011101110111",
				"100010001000",
				"100110011001",
				"100110011001",
				"101010101010",
				"101010101010",
				"100110011001",
				"100110011010",
				"101010101011",
				"101010111011",
				"101010111100",
				"101010111011",
				"101010111100",
				"101010111100",
				"100110101010",
				"011110011010",
				"101011001101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"101111011110",
				"110011011111",
				"101010111100",
				"100010001010",
				"101110111100",
				"111011101111",
				"101111001101",
				"101010111101",
				"101011001110",
				"101011011110",
				"100111011110",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101111101111",
				"110011101111",
				"101110111101",
				"011110001010",
				"101011011110",
				"100011011110",
				"100011011110",
				"100111011111",
				"100111101111",
				"101011011111",
				"101011101111",
				"101011101111",
				"101111101111",
				"101011011111",
				"100111011110",
				"101011011110",
				"110011101111",
				"110011101111",
				"101111011111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111101111",
				"101111101110",
				"110011011110",
				"101110111100",
				"011001010111",
				"011001010111",
				"100010001010",
				"101111011110",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011111",
				"101011101111",
				"101011001110",
				"011001111001",
				"010001010110",
				"011110011010",
				"011110011010",
				"100010101100",
				"100010101100",
				"011110011100",
				"011010001011",
				"011010011011",
				"011110111101",
				"011010101100",
				"011010101100",
				"011110111101",
				"100011001110",
				"100011001111",
				"011111001110",
				"011111001110",
				"100011011111",
				"011111001110",
				"011111001110",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"101011011111",
				"101011101111",
				"100011011110",
				"011010111100",
				"011010111101",
				"011111001110",
				"011111001101",
				"011111001110",
				"011111001110",
				"011111001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001110",
				"100011001110",
				"100011001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011110111101",
				"011110111100",
				"011110111100",
				"011110011010",
				"010001010111",
				"001101000110",
				"011001101000",
				"011110001010",
				"011110011011",
				"100011001101",
				"010110101100",
				"011011001110",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011010111100",
				"011010111100",
				"011010111100",
				"011111001100",
				"011110111100",
				"100011001100",
				"100111001101",
				"011010001001",
				"010001100111",
				"011010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101100",
				"011110101100",
				"011110101100",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111100",
				"011010111011",
				"011010111011",
				"011010111011",
				"011110111100",
				"011010101011",
				"010110011010",
				"011010101010",
				"011110101011",
				"011010011011",
				"011010011011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010101011",
				"010110101011",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110101011",
				"011010111011",
				"011010111011",
				"010110101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110101011",
				"010010001001",
				"010010011010",
				"010010011010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"011110111011",
				"100010111100",
				"011010011010",
				"011010011001",
				"100010101011",
				"100010011010",
				"011001111000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100000000",
				"000100010001",
				"001000010001",
				"001100100010",
				"010000110011",
				"010001000100",
				"010101000100",
				"010101010100",
				"010101010101",
				"011001100101",
				"010101010101",
				"011101110110",
				"011110000111",
				"100010001000",
				"100110011001",
				"101010101010",
				"100110011010",
				"100010011001",
				"100110011010",
				"101010111011",
				"101010101011",
				"101010111011",
				"101110111100",
				"101010111100",
				"100110101011",
				"011110001001",
				"100110111011",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011001110",
				"101111001110",
				"110011011110",
				"110011001110",
				"100010001001",
				"011001101000",
				"101010101011",
				"101110111101",
				"101010111100",
				"101011001101",
				"101011011110",
				"100111011111",
				"100111011111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101110",
				"101011011110",
				"101111101111",
				"110011011111",
				"011110001010",
				"100010111100",
				"100111011110",
				"100111011110",
				"100011011110",
				"100111011111",
				"101011011111",
				"101011011111",
				"101111011111",
				"101111011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101111101111",
				"110011101111",
				"110011101111",
				"101111101111",
				"101111101111",
				"110011111111",
				"110011111111",
				"110011101110",
				"101111011101",
				"100010001001",
				"011001010110",
				"011101100111",
				"100110101011",
				"101111011110",
				"101011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"100111011111",
				"101111011111",
				"100010011010",
				"010101010111",
				"011001111000",
				"011001111000",
				"011001111001",
				"011110001011",
				"011110001100",
				"100010101101",
				"100010111101",
				"100011001110",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111001111",
				"011111001110",
				"011111001110",
				"011011001110",
				"011111001110",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100111011111",
				"100111101111",
				"100011001110",
				"011111001101",
				"011111001101",
				"011111001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"100011001110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011011110",
				"100011011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011001110",
				"100011001101",
				"011110111100",
				"011110101100",
				"011010101100",
				"011010101011",
				"011110101011",
				"100110111100",
				"100010011010",
				"011001101000",
				"010101101000",
				"011010001010",
				"011110011011",
				"100011001101",
				"010110101100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011111001101",
				"011111001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001100",
				"011110111100",
				"011110111100",
				"011010111100",
				"011010111011",
				"011110111011",
				"100010101011",
				"100010101011",
				"011110001010",
				"010101111000",
				"010110011010",
				"011010101011",
				"011010111100",
				"011010101100",
				"011110111100",
				"011010111100",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"011010111011",
				"011010111100",
				"011010111011",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"011010111011",
				"011110111100",
				"011010101011",
				"011010111011",
				"011110111100",
				"011010101010",
				"011010011010",
				"011110101011",
				"100010111100",
				"011110101011",
				"011110101100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101100",
				"011010101011",
				"010110011010",
				"010010011010",
				"010010011010",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010111011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111100",
				"011010101011",
				"011010101011",
				"011010111011",
				"011111001100",
				"011010101011",
				"010010001001",
				"001110001001",
				"010010011010",
				"010110101011",
				"010110011010",
				"010110101011",
				"011010111100",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010111011",
				"011010101011",
				"011010101011",
				"010110011001",
				"010110001001",
				"011110101011",
				"100010111011",
				"100010101011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000010001",
				"001000100010",
				"001100110011",
				"010000110011",
				"010001000100",
				"010001000100",
				"010101010100",
				"011001100110",
				"011101110110",
				"100010000111",
				"100110011001",
				"101010101010",
				"100110011001",
				"100010011001",
				"100110101010",
				"101010101011",
				"101010111011",
				"101010101011",
				"101010111011",
				"101010111011",
				"100010011001",
				"100010011010",
				"101010111100",
				"101111011101",
				"101011001101",
				"101011011110",
				"101011011110",
				"101011001110",
				"101011001110",
				"101111001101",
				"110111011110",
				"101010101100",
				"010001000110",
				"011001101000",
				"101111001101",
				"101011001101",
				"101011001101",
				"101011011110",
				"101011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"101011101111",
				"101011101110",
				"101011011110",
				"101111011110",
				"110111101111",
				"100110101100",
				"011110011011",
				"100111001110",
				"100111011110",
				"100011001110",
				"100111011110",
				"101011011110",
				"101011011111",
				"101111011111",
				"101111011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101111011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101111",
				"110011101110",
				"101111001100",
				"011001100111",
				"010101000101",
				"100001111001",
				"101110111101",
				"101111011111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100011011111",
				"100011101111",
				"100011101111",
				"100011011111",
				"100011001110",
				"101011011110",
				"101111001101",
				"100010001001",
				"100010001001",
				"100010001001",
				"100010001010",
				"100110011100",
				"101010111110",
				"101111001111",
				"101011011111",
				"100011001111",
				"100011001111",
				"011111001111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111001110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011011001110",
				"011111011110",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100111101111",
				"100111101111",
				"011111001101",
				"011110111101",
				"100011001110",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"011111011101",
				"011111011110",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011001110",
				"100011001110",
				"011110111100",
				"011110111100",
				"011010101100",
				"011010101011",
				"011010101100",
				"011110111100",
				"011111001101",
				"100011001101",
				"100110111101",
				"101111011110",
				"100110111100",
				"010101111000",
				"010101111001",
				"011110011011",
				"011110111101",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110101011",
				"100010101011",
				"100110101011",
				"100010011010",
				"010101101000",
				"010010001001",
				"011010101011",
				"011010111100",
				"011010101100",
				"011110111101",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010101011",
				"011010111100",
				"011110111100",
				"011010101011",
				"011010011010",
				"011110011010",
				"100010101011",
				"100010101100",
				"100010111100",
				"011110111100",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010010001001",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010111011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"011010101011",
				"011010101011",
				"011110111100",
				"010110011010",
				"001110001001",
				"010010001001",
				"010110011010",
				"010110011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101100",
				"011010111100",
				"011010111100",
				"011010101011",
				"011010111100",
				"010010011010",
				"010110011010",
				"011010011010",
				"010110011010",
				"010110011001",
				"011010011010",
				"100010111011",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010000",
				"000100010001",
				"001000100001",
				"001000100010",
				"001000100010",
				"001101000011",
				"010001010100",
				"010101010101",
				"011101110111",
				"100110011001",
				"100010001000",
				"100010011001",
				"100110101010",
				"101010101011",
				"101010101010",
				"100110011010",
				"101010111011",
				"101110111100",
				"100110101011",
				"011110001001",
				"100110111100",
				"101111001101",
				"101011001101",
				"101011001101",
				"101111011110",
				"101111001110",
				"101011001101",
				"101111001101",
				"110011001101",
				"110011001101",
				"011001100111",
				"011001100111",
				"101111001101",
				"101010111101",
				"101111011111",
				"101011011110",
				"100111011111",
				"100111011111",
				"100111011111",
				"100111101111",
				"101011101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"110011101111",
				"101111011111",
				"011110011011",
				"100111001101",
				"100111011110",
				"100111001110",
				"100111011110",
				"101011011110",
				"101011011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101011011110",
				"101011011110",
				"110011101111",
				"110111101111",
				"110011101111",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101110",
				"110011101110",
				"110111111111",
				"011001111000",
				"010101010110",
				"100010001010",
				"101111001110",
				"101011011110",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111101111",
				"100011101111",
				"100011101111",
				"100011101111",
				"100011011110",
				"101011011110",
				"110011001101",
				"100010001000",
				"011001010110",
				"011101111000",
				"100010001011",
				"100110101101",
				"101010111110",
				"100111001111",
				"100011001111",
				"011111001110",
				"011111001111",
				"011111001111",
				"011111001110",
				"011011001110",
				"011011001110",
				"011111001110",
				"011111011111",
				"011111011111",
				"011111001110",
				"011111001110",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"011111011111",
				"011111011110",
				"100011101111",
				"011111011110",
				"100011011110",
				"100111101111",
				"100011001110",
				"011110111100",
				"100111001110",
				"100111001101",
				"100111001101",
				"100111001101",
				"100011001101",
				"100011001101",
				"100011001101",
				"100011011110",
				"100011011110",
				"100011011110",
				"100111011110",
				"100111011111",
				"100111011111",
				"100111011110",
				"100011001101",
				"011110111100",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010111100",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111001101",
				"100011001101",
				"100011001101",
				"100111001101",
				"101011011110",
				"011110101100",
				"010101111001",
				"010110001001",
				"011110111100",
				"011110111101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011010111100",
				"011110111100",
				"011110111011",
				"011110101011",
				"100110111100",
				"100010101011",
				"011001111001",
				"010101111000",
				"010110011010",
				"011010111100",
				"011010111100",
				"011010101100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011011001100",
				"011011001100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"011010111100",
				"011010111011",
				"010110101011",
				"011110111011",
				"011110011010",
				"010101111000",
				"010001010111",
				"011001111001",
				"011010001001",
				"010110001001",
				"010010001001",
				"010010001001",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110011010",
				"010110101011",
				"011010101011",
				"010110011010",
				"011110111100",
				"011010101011",
				"010110011010",
				"010010001001",
				"010110001010",
				"011010101011",
				"011010101011",
				"010110011010",
				"011010011011",
				"011010101011",
				"011010101011",
				"011110111100",
				"011110111100",
				"011110111100",
				"011010101100",
				"010110101011",
				"010010011010",
				"010010001001",
				"010110011011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"000100100001",
				"001000100010",
				"010001000100",
				"011001100110",
				"100010001000",
				"100010011001",
				"100110101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010101010",
				"101010111011",
				"101010111011",
				"011110001001",
				"100010011010",
				"101010111100",
				"101111001101",
				"101011001101",
				"101111001110",
				"101111011110",
				"101111001101",
				"101111001101",
				"101111001101",
				"110011011110",
				"100110101010",
				"011001100111",
				"100110101011",
				"110011011110",
				"101111011110",
				"101011011110",
				"100111011110",
				"100111011111",
				"100111011111",
				"101011101111",
				"101011101111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101111101111",
				"101111011111",
				"110111101111",
				"100110111100",
				"100110111101",
				"101111011111",
				"100111001101",
				"101011011110",
				"101011011110",
				"101111011111",
				"101111011111",
				"101111011111",
				"110011101111",
				"101111101111",
				"101111101111",
				"101111011110",
				"110011011111",
				"101111011110",
				"101011001101",
				"101011001101",
				"101011001110",
				"101111011110",
				"110011101111",
				"111011111111",
				"110111101111",
				"010101010111",
				"011110001001",
				"101111001110",
				"100111001110",
				"100011011110",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100011101111",
				"100011101111",
				"100111011110",
				"101011011110",
				"110011011110",
				"101010011010",
				"011001010110",
				"011101111000",
				"100010001010",
				"100110101101",
				"101011001111",
				"100111001111",
				"011110111110",
				"011111001110",
				"011111001111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111001111",
				"011111011111",
				"011111011111",
				"011111011110",
				"100011011111",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011111",
				"011111011111",
				"011111011111",
				"011111011111",
				"011111011110",
				"011111011110",
				"100011011111",
				"100011011110",
				"100011011110",
				"100111011110",
				"100010111101",
				"100010111100",
				"101011001110",
				"101111011110",
				"101011001110",
				"101011001110",
				"100111001110",
				"100111011110",
				"100111011111",
				"100111011110",
				"100111011110",
				"100011001110",
				"100011001101",
				"011110111100",
				"010110011011",
				"010110011010",
				"010110011010",
				"010110011011",
				"011010111100",
				"011110111101",
				"011111001101",
				"011111011110",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111011101",
				"100011011110",
				"100011001101",
				"100111011110",
				"100111011110",
				"100010111101",
				"011010101011",
				"010110011010",
				"011110101100",
				"011110111101",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011110111100",
				"011110111100",
				"100011001101",
				"100011001101",
				"100010111100",
				"100010101011",
				"011110001001",
				"011001111000",
				"010001100111",
				"010110011010",
				"011010101011",
				"010110101011",
				"011010111100",
				"011110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"011010111011",
				"011010101011",
				"011110101011",
				"011001111001",
				"001101000110",
				"010101101000",
				"011010001001",
				"011010011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110011010",
				"010110101011",
				"011010101011",
				"011010101011",
				"011110101011",
				"011010101011",
				"010110011010",
				"011010011010",
				"011010011011",
				"011010011011",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110101100",
				"011110111100",
				"011010101100",
				"010110011011",
				"010010001010",
				"010010001001",
				"010110011011",
				"010110011010",
				"010110101011",
				"010110011011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000100010001",
				"001000100010",
				"001100110011",
				"011001100110",
				"100010001000",
				"100110011001",
				"101010101010",
				"101010011010",
				"101010011010",
				"101010101011",
				"101010101011",
				"100110011010",
				"100010011010",
				"100110111011",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111001110",
				"101011001101",
				"101111001101",
				"101011001101",
				"110011011110",
				"101010111100",
				"011101111000",
				"100010011010",
				"101111001101",
				"101011001101",
				"101011011110",
				"100111011110",
				"100111011111",
				"100111011111",
				"101011011111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101011011110",
				"110011101111",
				"101010111101",
				"100110101100",
				"101111011111",
				"101011011110",
				"101011011110",
				"101011011110",
				"101111011111",
				"110011011111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101111101111",
				"100111001101",
				"101011001110",
				"101111001110",
				"101011001110",
				"101111011110",
				"101111011110",
				"101111011110",
				"101111101111",
				"110111101111",
				"110111101111",
				"011101111001",
				"011110001010",
				"101011001110",
				"100111001110",
				"100011011111",
				"100011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100011101111",
				"100011101111",
				"100011011110",
				"101011011101",
				"110011011101",
				"101010011010",
				"011001010110",
				"011101111000",
				"100010011011",
				"100110111101",
				"101011001111",
				"100111001111",
				"011111001111",
				"011111011111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"100011011111",
				"100011011111",
				"100011011111",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011111",
				"011111011111",
				"100011011111",
				"100011011110",
				"100011001110",
				"100111001110",
				"100010111100",
				"011110011011",
				"100010011011",
				"100110111100",
				"101010111101",
				"101011001110",
				"101011001110",
				"100010111101",
				"011110111100",
				"011010101011",
				"011010101011",
				"010110011011",
				"010110011011",
				"011010011011",
				"010110011011",
				"011010101100",
				"011110111101",
				"100011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011011001101",
				"011011011101",
				"011111011110",
				"011111011110",
				"011011001101",
				"011111011101",
				"100011011110",
				"100011001110",
				"100011001101",
				"011110101100",
				"011010101011",
				"011110111101",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001100",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111101",
				"011110111101",
				"011110111100",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010011010",
				"010101100111",
				"010001010111",
				"010101100111",
				"010101111000",
				"010110011010",
				"010110101011",
				"010110101011",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110111011",
				"010110101011",
				"011010101011",
				"011110101011",
				"011110011010",
				"011001111000",
				"010101101000",
				"011010001001",
				"011010011010",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"010110101011",
				"011010101011",
				"010110011010",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010011010",
				"011010011010",
				"011010011011",
				"011110101100",
				"011010011011",
				"011010011010",
				"010110001001",
				"010010001001",
				"010010001001",
				"010010001010",
				"010110011010",
				"010110011011",
				"010110011011",
				"010110011011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010110011010",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"000000000000",
				"001100110011",
				"011001100110",
				"100010001000",
				"101010101010",
				"101010011010",
				"100110011001",
				"101010101010",
				"101010101010",
				"101010101011",
				"100010011010",
				"100110101011",
				"101011001100",
				"101011001101",
				"101011001101",
				"101111001110",
				"101011001101",
				"101011001101",
				"101011001101",
				"101111011101",
				"101111011101",
				"100010011001",
				"011110001001",
				"101010111100",
				"101011001101",
				"101011011110",
				"100111011110",
				"100111011110",
				"100111011111",
				"101011011111",
				"101011011111",
				"101011011110",
				"101011011110",
				"101011011111",
				"101011011110",
				"101011011110",
				"110011101111",
				"110011011110",
				"100110101100",
				"101111011110",
				"101111101111",
				"101011011111",
				"101011011110",
				"110011101111",
				"110011101111",
				"110011101111",
				"101111011111",
				"101011001101",
				"100111001101",
				"100111001101",
				"101011001110",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011111",
				"101111011110",
				"101111011110",
				"110011011111",
				"110111101111",
				"100110011011",
				"011001111001",
				"100110111110",
				"100111001110",
				"100011011111",
				"100011011111",
				"100111101111",
				"100111101111",
				"100111101111",
				"100111101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"101011101111",
				"100111101111",
				"100111101111",
				"100111011111",
				"100111011111",
				"100111011111",
				"100011101111",
				"011111101111",
				"100011011110",
				"101011011101",
				"110011011101",
				"101010011010",
				"011001010110",
				"011001111000",
				"100010011011",
				"100111001110",
				"100111001111",
				"100011011111",
				"100011011111",
				"100011101111",
				"100011011111",
				"100011101111",
				"100111101111",
				"100011101111",
				"100011011111",
				"100011011111",
				"100011011111",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"100011011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"011111011110",
				"100011101111",
				"011111001110",
				"100011001110",
				"100111011110",
				"100111001110",
				"101011001101",
				"011110001010",
				"010101100111",
				"011001111000",
				"011001111001",
				"011001111001",
				"011010001010",
				"011010011010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011011",
				"011010101100",
				"011110111101",
				"011110111101",
				"011111001101",
				"100011001110",
				"100011001110",
				"011111011110",
				"011111011110",
				"011111001110",
				"011011001101",
				"011011001101",
				"011011011101",
				"011011011110",
				"011011011110",
				"011011011101",
				"011011011101",
				"011011011101",
				"011111011101",
				"100011011110",
				"100111011110",
				"100010111100",
				"011010011011",
				"011110111101",
				"011010111100",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011011001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011011001101",
				"011010111100",
				"011010111100",
				"011110111101",
				"011110111101",
				"011110111101",
				"011111001101",
				"011111001101",
				"011111001101",
				"011110111100",
				"011010101011",
				"011010101011",
				"010110001001",
				"001101010110",
				"010001000110",
				"010101100111",
				"010101111000",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"011010111100",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110111100",
				"010110111011",
				"010110111011",
				"010110101011",
				"011010101010",
				"011110101011",
				"100010011011",
				"011110001001",
				"011001111000",
				"011010001001",
				"011010011010",
				"010110011010",
				"011010101011",
				"011010111011",
				"011010101100",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"011010101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101010",
				"010110101010",
				"011010101011",
				"011010101011",
				"011010101011",
				"011010011011",
				"011110101011",
				"011010011011",
				"010001111000",
				"001101010111",
				"010001101000",
				"010001111000",
				"010001111000",
				"010001111000",
				"010001111001",
				"010110001010",
				"010110011010",
				"010110001010",
				"010110001010",
				"010110011010",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110101011",
				"010110011010",
				"010110011010",
				"010110011010",
				"010010011010",
				"1111111111111");  -- bits de test

BEGIN
    PROCESS(RST, IS_SERPENT, XMAX, YMAX, HCOUNT, VCOUNT)
    BEGIN
        IF (RST = '1') THEN
            RED <= (OTHERS => '0');
            GREEN <= (OTHERS => '0');
            BLUE <= (OTHERS => '0');
            DEP_IMA <= '0';
        ELSE 
            IF (IS_SERPENT = '1') THEN
				IF (HCOUNT = XMAX AND VCOUNT = YMAX) THEN
					IF (data_vector(HCOUNT * VCOUNT) = data_vector(189000)) THEN
						DEP_IMA <= '0';    -- Si la dernière valeur est la même que la valeur actuelle
					ELSE
						DEP_IMA <= '1';    -- Si la dernière valeur est différente de la valeur actuelle
					END IF;
                ELSIF (HCOUNT * VCOUNT < 189000) THEN
                    RED <= data_vector(HCOUNT * VCOUNT)(0 DOWNTO 3);
                    GREEN <= data_vector(HCOUNT * VCOUNT)(4 DOWNTO 6);
                    BLUE <= data_vector(HCOUNT * VCOUNT)(7 DOWNTO 11);
                END IF;
            END IF;
        END IF;
    END PROCESS;
END rtl;
